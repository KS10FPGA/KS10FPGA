////////////////////////////////////////////////////////////////////
//!
//! KS-10 Processor
//!
//! \brief
//!      Dispatch ROM (DROM)
//!
//! \details
//!
//! \todo
//!
//! \file
//!      drom.v
//!
//! \author
//!      Rob Doyle - doyle (at) cox (dot) net
//!
////////////////////////////////////////////////////////////////////
//
//  Copyright (C) 2009, 2012 Rob Doyle
//
// This source file may be used and distributed without
// restriction provided that this copyright statement is not
// removed from the file and that any derivative work contains
// the original copyright notice and the associated disclaimer.
//
// This source file is free software; you can redistribute it
// and/or modify it under the terms of the GNU Lesser General
// Public License as published by the Free Software Foundation;
// version 2.1 of the License.
//
// This source is distributed in the hope that it will be
// useful, but WITHOUT ANY WARRANTY; without even the implied
// warranty of MERCHANTABILITY or FITNESS FOR A PARTICULAR
// PURPOSE. See the GNU Lesser General Public License for more
// details.
//
// You should have received a copy of the GNU Lesser General
// Public License along with this source; if not, download it
// from http://www.gnu.org/licenses/lgpl.txt
//
////////////////////////////////////////////////////////////////////
//
// Comments are formatted for doxygen
//

`include "crom.vh"
`include "drom.vh"

module DROM(clk, rst, clken, dbus, crom, drom);

   parameter  cromWidth = `CROM_WIDTH;
   parameter  dromWidth = `DROM_WIDTH;

   input                      clk;      // Clock
   input                      rst;      // Reset
   input                      clken;    // Clock Enable
   input      [0:35]          dbus;     // DBUS
   input      [0:cromWidth-1] crom;     // Control ROM
   output reg [0:dromWidth-1] drom;     // Dispatch ROM Output

   //
   // The DROM in the KS10 is asynchronous.  That won't work in an FPGA
   // implementation.  Fortunately the DROM is addressed by the Instruction
   // Register (IR) which is synchronous.  Therefore when we load the IR
   // we also load the address of the DROM.
   //
   
   wire loadIR = `cromSPEC_EN_40 & (`cromSPEC_SEL == `cromSPEC_SEL_LOADIR);
   wire [0:8] addr = dbus[0:8];

   //
   // Dispatch ROM (DROM)
   //  DPEA/E98
   //  DPEA/E117
   //  DPEA/E110
   //

   reg [0:dromWidth-1] DROM[0:511];
   
   initial
     begin
        DROM[  0] = 36'o0000_1556_2100;
        DROM[  1] = 36'o0001_1740_2100;
        DROM[  2] = 36'o0002_1740_2100;
        DROM[  3] = 36'o0003_1740_2100;
        DROM[  4] = 36'o0002_1741_2100;
        DROM[  5] = 36'o0005_1740_2100;
        DROM[  6] = 36'o0006_1740_2100;
        DROM[  7] = 36'o0007_1740_2100;
        DROM[  8] = 36'o0001_1742_2100;
        DROM[  9] = 36'o0004_1742_2100;
        DROM[ 10] = 36'o0001_1743_2100;
        DROM[ 11] = 36'o0000_1743_2100;
        DROM[ 12] = 36'o0001_1744_2100;
        DROM[ 13] = 36'o0000_1744_2100;
        DROM[ 14] = 36'o0002_1744_2100;
        DROM[ 15] = 36'o0003_1744_2100;
        DROM[ 16] = 36'o0000_1746_2100;
        DROM[ 17] = 36'o0000_1747_2100;
        DROM[ 18] = 36'o0000_1750_2100;
        DROM[ 19] = 36'o0000_1751_2100;
        DROM[ 20] = 36'o0001_1751_2100;
        DROM[ 21] = 36'o0002_1751_2100;
        DROM[ 22] = 36'o0004_1751_2100;
        DROM[ 23] = 36'o0010_1751_2100;
        DROM[ 24] = 36'o0000_1557_2100;
        DROM[ 25] = 36'o0001_1557_2100;
        DROM[ 26] = 36'o0002_1557_2100;
        DROM[ 27] = 36'o0003_1557_2100;
        DROM[ 28] = 36'o0004_1557_2100;
        DROM[ 29] = 36'o0005_1557_2100;
        DROM[ 30] = 36'o0006_1557_2100;
        DROM[ 31] = 36'o0007_1557_2100;
        DROM[ 32] = 36'o0000_1556_2100;
        DROM[ 33] = 36'o0000_1556_2100;
        DROM[ 34] = 36'o0000_1556_2100;
        DROM[ 35] = 36'o0000_1556_2100;
        DROM[ 36] = 36'o0000_1556_2100;
        DROM[ 37] = 36'o0000_1556_2100;
        DROM[ 38] = 36'o0000_1556_2100;
        DROM[ 39] = 36'o0000_1556_2100;
        DROM[ 40] = 36'o0000_1556_2100;
        DROM[ 41] = 36'o0000_1556_2100;
        DROM[ 42] = 36'o0000_1556_2100;
        DROM[ 43] = 36'o0000_1556_2100;
        DROM[ 44] = 36'o0000_1556_2100;
        DROM[ 45] = 36'o0000_1556_2100;
        DROM[ 46] = 36'o0000_1556_2100;
        DROM[ 47] = 36'o0000_1556_2100;
        DROM[ 48] = 36'o0000_1556_2100;
        DROM[ 49] = 36'o0000_1556_2100;
        DROM[ 50] = 36'o0000_1556_2100;
        DROM[ 51] = 36'o0000_1556_2100;
        DROM[ 52] = 36'o0000_1556_2100;
        DROM[ 53] = 36'o0000_1556_2100;
        DROM[ 54] = 36'o0000_1556_2100;
        DROM[ 55] = 36'o0000_1556_2100;
        DROM[ 56] = 36'o0000_1556_2100;
        DROM[ 57] = 36'o0000_1556_2100;
        DROM[ 58] = 36'o0000_1556_2100;
        DROM[ 59] = 36'o0000_1556_2100;
        DROM[ 60] = 36'o0000_1556_2100;
        DROM[ 61] = 36'o0000_1556_2100;
        DROM[ 62] = 36'o0000_1556_2100;
        DROM[ 63] = 36'o0000_1556_2100;
        DROM[ 64] = 36'o0000_1556_2100;
        DROM[ 65] = 36'o0000_1661_2100;
        DROM[ 66] = 36'o0000_1662_2100;
        DROM[ 67] = 36'o0000_1663_2100;
        DROM[ 68] = 36'o0000_1664_2100;
        DROM[ 69] = 36'o0000_1551_3000;
        DROM[ 70] = 36'o0000_1666_2100;
        DROM[ 71] = 36'o0000_1667_2100;
        DROM[ 72] = 36'o1100_1637_1100;
        DROM[ 73] = 36'o1100_1635_1100;
        DROM[ 74] = 36'o1105_1631_1100;
        DROM[ 75] = 36'o1105_1636_1100;
        DROM[ 76] = 36'o0205_1457_1100;
        DROM[ 77] = 36'o0205_1615_1100;
        DROM[ 78] = 36'o0205_1566_1100;
        DROM[ 79] = 36'o0205_1627_1100;
        DROM[ 80] = 36'o0205_1505_1100;
        DROM[ 81] = 36'o0215_1434_1100;
        DROM[ 82] = 36'o0701_1626_1100;
        DROM[ 83] = 36'o0000_1467_3100;
        DROM[ 84] = 36'o0300_1567_0100;
        DROM[ 85] = 36'o0100_1565_0500;
        DROM[ 86] = 36'o0711_1626_1100;
        DROM[ 87] = 36'o0011_1616_1100;
        DROM[ 88] = 36'o0000_1660_2100;
        DROM[ 89] = 36'o0001_1660_2100;
        DROM[ 90] = 36'o0001_1621_2100;
        DROM[ 91] = 36'o0015_1610_1100;
        DROM[ 92] = 36'o0000_1620_1500;
        DROM[ 93] = 36'o0000_1624_1100;
        DROM[ 94] = 36'o0000_1630_1500;
        DROM[ 95] = 36'o0000_1634_1100;
        DROM[ 96] = 36'o0701_1577_1100;
        DROM[ 97] = 36'o0002_1660_2100;
        DROM[ 98] = 36'o0702_1577_1700;
        DROM[ 99] = 36'o0703_1577_1700;
        DROM[100] = 36'o0711_1577_1100;
        DROM[101] = 36'o0611_1577_0100;
        DROM[102] = 36'o0712_1577_1700;
        DROM[103] = 36'o0713_1577_1700;
        DROM[104] = 36'o0701_1576_1100;
        DROM[105] = 36'o0003_1660_2100;
        DROM[106] = 36'o0702_1576_1700;
        DROM[107] = 36'o0703_1576_1700;
        DROM[108] = 36'o0711_1576_1100;
        DROM[109] = 36'o0611_1576_0100;
        DROM[110] = 36'o0712_1576_1700;
        DROM[111] = 36'o0713_1576_1700;
        DROM[112] = 36'o0701_1570_1100;
        DROM[113] = 36'o0004_1660_2100;
        DROM[114] = 36'o0702_1570_1700;
        DROM[115] = 36'o0703_1570_1700;
        DROM[116] = 36'o0711_1570_1100;
        DROM[117] = 36'o0611_1570_0100;
        DROM[118] = 36'o0712_1570_1700;
        DROM[119] = 36'o0713_1570_1700;
        DROM[120] = 36'o0701_1574_1100;
        DROM[121] = 36'o0005_1660_2100;
        DROM[122] = 36'o0702_1574_1700;
        DROM[123] = 36'o0703_1574_1700;
        DROM[124] = 36'o0711_1574_1100;
        DROM[125] = 36'o0611_1574_0100;
        DROM[126] = 36'o0712_1574_1700;
        DROM[127] = 36'o0713_1574_1700;
        DROM[128] = 36'o1015_1515_1100;
        DROM[129] = 36'o0015_1515_3000;
        DROM[130] = 36'o0116_1404_0700;
        DROM[131] = 36'o0004_1504_1700;
        DROM[132] = 36'o1015_1402_1100;
        DROM[133] = 36'o0015_1402_3000;
        DROM[134] = 36'o0116_1402_0700;
        DROM[135] = 36'o0004_1402_1700;
        DROM[136] = 36'o1015_1405_1100;
        DROM[137] = 36'o0015_1405_3000;
        DROM[138] = 36'o0116_1405_0700;
        DROM[139] = 36'o0004_1405_1700;
        DROM[140] = 36'o1015_1403_1100;
        DROM[141] = 36'o0015_1515_3000;
        DROM[142] = 36'o0116_1403_0700;
        DROM[143] = 36'o0004_1403_1700;
        DROM[144] = 36'o1015_1641_1100;
        DROM[145] = 36'o0015_1641_3000;
        DROM[146] = 36'o0016_1641_1700;
        DROM[147] = 36'o0017_1641_1700;
        DROM[148] = 36'o1005_1571_1100;
        DROM[149] = 36'o0005_1571_3000;
        DROM[150] = 36'o0016_1571_1700;
        DROM[151] = 36'o0006_1571_1700;
        DROM[152] = 36'o1005_1600_1100;
        DROM[153] = 36'o0005_1600_3000;
        DROM[154] = 36'o0016_1600_1700;
        DROM[155] = 36'o0006_1600_1700;
        DROM[156] = 36'o1005_1601_1100;
        DROM[157] = 36'o0005_1601_3000;
        DROM[158] = 36'o0016_1601_1700;
        DROM[159] = 36'o0006_1601_1700;
        DROM[160] = 36'o0400_1622_1000;
        DROM[161] = 36'o0400_1632_1000;
        DROM[162] = 36'o0400_1612_1000;
        DROM[163] = 36'o0000_1462_2100;
        DROM[164] = 36'o0000_1466_3000;
        DROM[165] = 36'o0500_1470_1000;
        DROM[166] = 36'o0500_1464_1000;
        DROM[167] = 36'o0000_1665_2100;
        DROM[168] = 36'o0015_1406_1500;
        DROM[169] = 36'o0000_1640_2100;
        DROM[170] = 36'o0005_1547_2100;
        DROM[171] = 36'o0001_1547_2100;
        DROM[172] = 36'o0000_1520_6000;
        DROM[173] = 36'o0000_1540_2100;
        DROM[174] = 36'o0000_1541_1100;
        DROM[175] = 36'o1215_1553_0100;
        DROM[176] = 36'o0000_1544_2100;
        DROM[177] = 36'o0002_1543_3100;
        DROM[178] = 36'o0002_1545_2100;
        DROM[179] = 36'o0000_1546_2100;
        DROM[180] = 36'o0000_1552_2100;
        DROM[181] = 36'o0000_1550_2100;
        DROM[182] = 36'o0000_1554_2100;
        DROM[183] = 36'o0000_1555_2100;
        DROM[184] = 36'o1015_1560_1100;
        DROM[185] = 36'o0015_1560_3000;
        DROM[186] = 36'o0016_1560_1700;
        DROM[187] = 36'o0017_1560_1700;
        DROM[188] = 36'o1015_1561_1100;
        DROM[189] = 36'o0015_1561_3000;
        DROM[190] = 36'o0016_1561_1700;
        DROM[191] = 36'o0017_1561_1700;
        DROM[192] = 36'o0000_1400_2100;
        DROM[193] = 36'o0001_1476_2100;
        DROM[194] = 36'o0002_1476_2100;
        DROM[195] = 36'o0003_1476_2100;
        DROM[196] = 36'o0004_1476_2100;
        DROM[197] = 36'o0005_1476_2100;
        DROM[198] = 36'o0006_1476_2100;
        DROM[199] = 36'o0007_1476_2100;
        DROM[200] = 36'o0000_1476_1100;
        DROM[201] = 36'o0001_1476_1100;
        DROM[202] = 36'o0002_1476_1100;
        DROM[203] = 36'o0003_1476_1100;
        DROM[204] = 36'o0004_1476_1100;
        DROM[205] = 36'o0005_1476_1100;
        DROM[206] = 36'o0006_1476_1100;
        DROM[207] = 36'o0007_1476_1100;
        DROM[208] = 36'o0000_1400_2100;
        DROM[209] = 36'o0001_1440_2100;
        DROM[210] = 36'o0002_1440_2100;
        DROM[211] = 36'o0003_1440_2100;
        DROM[212] = 36'o0004_1520_2100;
        DROM[213] = 36'o0005_1440_2100;
        DROM[214] = 36'o0006_1440_2100;
        DROM[215] = 36'o0007_1440_2100;
        DROM[216] = 36'o0000_1477_1100;
        DROM[217] = 36'o0001_1477_1100;
        DROM[218] = 36'o0002_1477_1100;
        DROM[219] = 36'o0003_1477_1100;
        DROM[220] = 36'o0004_1477_1100;
        DROM[221] = 36'o0005_1477_1100;
        DROM[222] = 36'o0006_1477_1100;
        DROM[223] = 36'o0007_1477_1100;
        DROM[224] = 36'o0000_1611_3000;
        DROM[225] = 36'o0001_1611_2100;
        DROM[226] = 36'o0002_1611_2100;
        DROM[227] = 36'o0003_1611_2100;
        DROM[228] = 36'o0004_1611_2100;
        DROM[229] = 36'o0005_1611_2100;
        DROM[230] = 36'o0006_1611_2100;
        DROM[231] = 36'o0007_1611_2100;
        DROM[232] = 36'o0000_1431_1500;
        DROM[233] = 36'o0001_1431_1500;
        DROM[234] = 36'o0002_1431_1500;
        DROM[235] = 36'o0003_1431_1500;
        DROM[236] = 36'o0004_1431_1500;
        DROM[237] = 36'o0005_1431_1500;
        DROM[238] = 36'o0006_1431_1500;
        DROM[239] = 36'o0007_1431_1500;
        DROM[240] = 36'o0000_1542_3000;
        DROM[241] = 36'o0001_1542_2100;
        DROM[242] = 36'o0002_1542_2100;
        DROM[243] = 36'o0003_1542_2100;
        DROM[244] = 36'o0004_1542_2100;
        DROM[245] = 36'o0005_1542_2100;
        DROM[246] = 36'o0006_1542_2100;
        DROM[247] = 36'o0007_1542_2100;
        DROM[248] = 36'o0000_1437_1500;
        DROM[249] = 36'o0001_1437_1500;
        DROM[250] = 36'o0002_1437_1500;
        DROM[251] = 36'o0003_1437_1500;
        DROM[252] = 36'o0004_1437_1500;
        DROM[253] = 36'o0005_1437_1500;
        DROM[254] = 36'o0006_1437_1500;
        DROM[255] = 36'o0007_1437_1500;
        DROM[256] = 36'o0015_1441_3000;
        DROM[257] = 36'o0015_1441_3000;
        DROM[258] = 36'o0016_1441_2700;
        DROM[259] = 36'o0017_1441_2700;
        DROM[260] = 36'o1015_1442_1100;
        DROM[261] = 36'o0015_1442_3000;
        DROM[262] = 36'o0016_1442_1700;
        DROM[263] = 36'o0017_1442_1700;
        DROM[264] = 36'o1015_1443_1100;
        DROM[265] = 36'o0015_1443_3000;
        DROM[266] = 36'o0016_1443_1700;
        DROM[267] = 36'o0017_1443_1700;
        DROM[268] = 36'o1015_1404_1100;
        DROM[269] = 36'o0015_1404_3000;
        DROM[270] = 36'o0016_1404_1700;
        DROM[271] = 36'o0017_1404_1700;
        DROM[272] = 36'o1015_1444_1100;
        DROM[273] = 36'o0015_1444_3000;
        DROM[274] = 36'o0016_1444_1700;
        DROM[275] = 36'o0017_1444_1700;
        DROM[276] = 36'o0000_1400_1100;
        DROM[277] = 36'o0000_1400_2100;
        DROM[278] = 36'o0116_1404_0700;
        DROM[279] = 36'o0116_1404_0700;
        DROM[280] = 36'o1015_1445_1100;
        DROM[281] = 36'o0015_1445_3000;
        DROM[282] = 36'o0016_1445_1700;
        DROM[283] = 36'o0017_1445_1700;
        DROM[284] = 36'o1015_1446_1100;
        DROM[285] = 36'o0015_1446_3000;
        DROM[286] = 36'o0016_1446_1700;
        DROM[287] = 36'o0017_1446_1700;
        DROM[288] = 36'o1015_1447_1100;
        DROM[289] = 36'o0015_1447_3000;
        DROM[290] = 36'o0016_1447_1700;
        DROM[291] = 36'o0017_1447_1700;
        DROM[292] = 36'o1015_1450_1100;
        DROM[293] = 36'o0015_1450_3000;
        DROM[294] = 36'o0016_1450_1700;
        DROM[295] = 36'o0017_1450_1700;
        DROM[296] = 36'o0015_1451_3000;
        DROM[297] = 36'o0015_1451_3000;
        DROM[298] = 36'o0016_1451_2700;
        DROM[299] = 36'o0017_1451_2700;
        DROM[300] = 36'o1015_1452_1100;
        DROM[301] = 36'o0015_1452_3000;
        DROM[302] = 36'o0016_1452_1700;
        DROM[303] = 36'o0017_1452_1700;
        DROM[304] = 36'o1015_1453_1100;
        DROM[305] = 36'o0015_1453_3000;
        DROM[306] = 36'o0016_1453_1700;
        DROM[307] = 36'o0017_1453_1700;
        DROM[308] = 36'o1015_1454_1100;
        DROM[309] = 36'o0015_1454_3000;
        DROM[310] = 36'o0016_1454_1700;
        DROM[311] = 36'o0017_1454_1700;
        DROM[312] = 36'o1015_1455_1100;
        DROM[313] = 36'o0015_1455_3000;
        DROM[314] = 36'o0016_1455_1700;
        DROM[315] = 36'o0017_1455_1700;
        DROM[316] = 36'o0015_1456_3000;
        DROM[317] = 36'o0015_1456_3000;
        DROM[318] = 36'o0016_1456_2700;
        DROM[319] = 36'o0017_1456_2700;
        DROM[320] = 36'o1015_1410_1100;
        DROM[321] = 36'o0015_1410_3000;
        DROM[322] = 36'o0016_1407_1700;
        DROM[323] = 36'o0004_1404_1700;
        DROM[324] = 36'o1015_1411_1100;
        DROM[325] = 36'o0015_1411_3000;
        DROM[326] = 36'o0016_1413_1700;
        DROM[327] = 36'o0004_1414_1700;
        DROM[328] = 36'o1015_1432_1100;
        DROM[329] = 36'o0015_1432_3000;
        DROM[330] = 36'o0116_1432_0700;
        DROM[331] = 36'o0004_1432_1700;
        DROM[332] = 36'o1015_1424_1100;
        DROM[333] = 36'o0015_1424_3000;
        DROM[334] = 36'o0116_1424_0700;
        DROM[335] = 36'o0004_1424_1700;
        DROM[336] = 36'o1015_1433_1100;
        DROM[337] = 36'o0015_1433_3000;
        DROM[338] = 36'o0116_1433_0700;
        DROM[339] = 36'o0004_1433_1700;
        DROM[340] = 36'o1015_1425_1100;
        DROM[341] = 36'o0015_1425_3000;
        DROM[342] = 36'o0116_1425_0700;
        DROM[343] = 36'o0004_1425_1700;
        DROM[344] = 36'o1015_1430_1100;
        DROM[345] = 36'o0015_1430_3000;
        DROM[346] = 36'o0116_1430_0700;
        DROM[347] = 36'o0004_1430_1700;
        DROM[348] = 36'o1015_1422_1100;
        DROM[349] = 36'o0015_1422_3000;
        DROM[350] = 36'o0116_1422_0700;
        DROM[351] = 36'o0004_1422_1700;
        DROM[352] = 36'o1015_1407_1100;
        DROM[353] = 36'o0015_1407_3000;
        DROM[354] = 36'o0016_1410_1700;
        DROM[355] = 36'o0004_1404_1700;
        DROM[356] = 36'o1015_1412_1100;
        DROM[357] = 36'o0015_1412_3000;
        DROM[358] = 36'o0016_1415_1700;
        DROM[359] = 36'o0004_1416_1700;
        DROM[360] = 36'o1015_1420_1100;
        DROM[361] = 36'o0015_1420_3000;
        DROM[362] = 36'o0116_1420_0700;
        DROM[363] = 36'o0004_1420_1700;
        DROM[364] = 36'o1015_1426_1100;
        DROM[365] = 36'o0015_1426_3000;
        DROM[366] = 36'o0116_1426_0700;
        DROM[367] = 36'o0004_1426_1700;
        DROM[368] = 36'o1015_1421_1100;
        DROM[369] = 36'o0015_1421_3000;
        DROM[370] = 36'o0116_1421_0700;
        DROM[371] = 36'o0004_1421_1700;
        DROM[372] = 36'o1015_1427_1100;
        DROM[373] = 36'o0015_1427_3000;
        DROM[374] = 36'o0116_1427_0700;
        DROM[375] = 36'o0004_1427_1700;
        DROM[376] = 36'o1015_1417_1100;
        DROM[377] = 36'o0015_1417_3000;
        DROM[378] = 36'o0116_1417_0700;
        DROM[379] = 36'o0004_1417_1700;
        DROM[380] = 36'o1015_1423_1100;
        DROM[381] = 36'o0015_1423_3000;
        DROM[382] = 36'o0116_1423_0700;
        DROM[383] = 36'o0004_1423_1700;
        DROM[384] = 36'o0000_1400_2100;
        DROM[385] = 36'o0000_1400_2100;
        DROM[386] = 36'o0000_1475_2100;
        DROM[387] = 36'o0000_1474_2100;
        DROM[388] = 36'o0000_1473_2100;
        DROM[389] = 36'o0000_1472_2100;
        DROM[390] = 36'o0004_1475_2100;
        DROM[391] = 36'o0004_1474_2100;
        DROM[392] = 36'o0000_1400_2100;
        DROM[393] = 36'o0000_1400_2100;
        DROM[394] = 36'o0000_1475_1100;
        DROM[395] = 36'o0000_1474_1100;
        DROM[396] = 36'o0000_1473_1100;
        DROM[397] = 36'o0000_1472_1100;
        DROM[398] = 36'o0004_1475_1100;
        DROM[399] = 36'o0004_1474_1100;
        DROM[400] = 36'o0005_1473_2100;
        DROM[401] = 36'o0005_1472_2100;
        DROM[402] = 36'o0001_1475_2100;
        DROM[403] = 36'o0001_1474_2100;
        DROM[404] = 36'o0001_1473_2100;
        DROM[405] = 36'o0001_1472_2100;
        DROM[406] = 36'o0005_1475_2100;
        DROM[407] = 36'o0005_1474_2100;
        DROM[408] = 36'o0005_1473_1100;
        DROM[409] = 36'o0005_1472_1100;
        DROM[410] = 36'o0001_1475_1100;
        DROM[411] = 36'o0001_1474_1100;
        DROM[412] = 36'o0001_1473_1100;
        DROM[413] = 36'o0001_1472_1100;
        DROM[414] = 36'o0005_1475_1100;
        DROM[415] = 36'o0005_1474_1100;
        DROM[416] = 36'o0006_1473_2100;
        DROM[417] = 36'o0006_1472_2100;
        DROM[418] = 36'o0002_1475_2100;
        DROM[419] = 36'o0002_1474_2100;
        DROM[420] = 36'o0002_1473_2100;
        DROM[421] = 36'o0002_1472_2100;
        DROM[422] = 36'o0006_1475_2100;
        DROM[423] = 36'o0006_1474_2100;
        DROM[424] = 36'o0006_1473_1100;
        DROM[425] = 36'o0006_1472_1100;
        DROM[426] = 36'o0002_1475_1100;
        DROM[427] = 36'o0002_1474_1100;
        DROM[428] = 36'o0002_1473_1100;
        DROM[429] = 36'o0002_1472_1100;
        DROM[430] = 36'o0006_1475_1100;
        DROM[431] = 36'o0006_1474_1100;
        DROM[432] = 36'o0007_1473_2100;
        DROM[433] = 36'o0007_1472_2100;
        DROM[434] = 36'o0003_1475_2100;
        DROM[435] = 36'o0003_1474_2100;
        DROM[436] = 36'o0003_1473_2100;
        DROM[437] = 36'o0003_1472_2100;
        DROM[438] = 36'o0007_1475_2100;
        DROM[439] = 36'o0007_1474_2100;
        DROM[440] = 36'o0007_1473_1100;
        DROM[441] = 36'o0007_1472_1100;
        DROM[442] = 36'o0003_1475_1100;
        DROM[443] = 36'o0003_1474_1100;
        DROM[444] = 36'o0003_1473_1100;
        DROM[445] = 36'o0003_1472_1100;
        DROM[446] = 36'o0007_1475_1100;
        DROM[447] = 36'o0007_1474_1100;
        DROM[448] = 36'o1200_1700_4100;
        DROM[449] = 36'o1200_1720_4100;
        DROM[450] = 36'o1216_1760_4700;
        DROM[451] = 36'o0003_1650_2100;
        DROM[452] = 36'o1200_1754_0100;
        DROM[453] = 36'o1200_1755_0100;
        DROM[454] = 36'o0006_1650_2100;
        DROM[455] = 36'o0007_1650_2100;
        DROM[456] = 36'o1210_1614_0100;
        DROM[457] = 36'o1214_1614_0100;
        DROM[458] = 36'o1210_1460_0100;
        DROM[459] = 36'o1210_1461_0100;
        DROM[460] = 36'o1210_1644_0100;
        DROM[461] = 36'o1214_1644_0100;
        DROM[462] = 36'o0006_1651_2100;
        DROM[463] = 36'o0007_1651_2100;
        DROM[464] = 36'o1200_1614_0100;
        DROM[465] = 36'o1204_1614_0100;
        DROM[466] = 36'o1200_1460_0100;
        DROM[467] = 36'o1200_1461_0100;
        DROM[468] = 36'o1200_1644_0100;
        DROM[469] = 36'o1204_1644_0100;
        DROM[470] = 36'o0006_1652_2100;
        DROM[471] = 36'o0007_1652_2100;
        DROM[472] = 36'o0000_1653_2100;
        DROM[473] = 36'o0001_1653_2100;
        DROM[474] = 36'o0002_1653_2100;
        DROM[475] = 36'o0003_1653_2100;
        DROM[476] = 36'o0004_1653_2100;
        DROM[477] = 36'o0005_1653_2100;
        DROM[478] = 36'o0006_1653_2100;
        DROM[479] = 36'o0007_1653_2100;
        DROM[480] = 36'o0000_1654_2100;
        DROM[481] = 36'o0001_1654_2100;
        DROM[482] = 36'o0002_1654_2100;
        DROM[483] = 36'o0003_1654_2100;
        DROM[484] = 36'o0004_1654_2100;
        DROM[485] = 36'o0005_1654_2100;
        DROM[486] = 36'o0006_1654_2100;
        DROM[487] = 36'o0007_1654_2100;
        DROM[488] = 36'o0000_1655_2100;
        DROM[489] = 36'o0001_1655_2100;
        DROM[490] = 36'o0002_1655_2100;
        DROM[491] = 36'o0003_1655_2100;
        DROM[492] = 36'o0004_1655_2100;
        DROM[493] = 36'o0005_1655_2100;
        DROM[494] = 36'o0006_1655_2100;
        DROM[495] = 36'o0007_1655_2100;
        DROM[496] = 36'o0000_1656_2100;
        DROM[497] = 36'o0001_1656_2100;
        DROM[498] = 36'o0002_1656_2100;
        DROM[499] = 36'o0003_1656_2100;
        DROM[500] = 36'o0004_1656_2100;
        DROM[501] = 36'o0005_1656_2100;
        DROM[502] = 36'o0006_1656_2100;
        DROM[503] = 36'o0007_1656_2100;
        DROM[504] = 36'o0000_1657_2100;
        DROM[505] = 36'o0001_1657_2100;
        DROM[506] = 36'o0002_1657_2100;
        DROM[507] = 36'o0003_1657_2100;
        DROM[508] = 36'o0004_1657_2100;
        DROM[509] = 36'o0005_1657_2100;
        DROM[510] = 36'o0006_1657_2100;
        DROM[511] = 36'o0007_1657_2100;
     end

   //
   // Synchronous ROM
   //

   always @(posedge clk)
     begin
        if (rst)
          drom <= 36'b0;
        else if (clken & loadIR)
          drom <= DROM[addr];
     end

endmodule
