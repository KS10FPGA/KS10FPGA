////////////////////////////////////////////////////////////////////////////////
//
// KS-10 Processor
//
// Brief
//   Debug Interface
//
// Details
//   This module provides KS10 breakpoint and instruction trace capabilities.
//   - the breakpoint is accomplished by examining the CPU Address Bus.
//   - the trace accesses the Program Counter (PC) and the Instruction Register
//     (IR).
//
// File
//   debug.v
//
// Author
//   Rob Doyle - doyle (at) cox (dot) net
//
////////////////////////////////////////////////////////////////////////////////
//
// Copyright (C) 2012-2017 Rob Doyle
//
// This source file may be used and distributed without restriction provided
// that this copyright statement is not removed from the file and that any
// derivative work contains the original copyright notice and the associated
// disclaimer.
//
// This source file is free software; you can redistribute it and/or modify it
// under the terms of the GNU Lesser General Public License as published by the
// Free Software Foundation; version 2.1 of the License.
//
// This source is distributed in the hope that it will be useful, but WITHOUT
// ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
// FITNESS FOR A PARTICULAR PURPOSE. See the GNU Lesser General Public License
// for more details.
//
// You should have received a copy of the GNU Lesser General Public License
// along with this source; if not, download it from
// http://www.gnu.org/licenses/lgpl.txt
//
////////////////////////////////////////////////////////////////////////////////

`default_nettype none
`timescale 1ns/1ps

module DEBUG (
      input  wire         rst,          // Reset
      input  wire         clk,          // Clock
      input  wire [ 0:35] cpuADDR,      // Backplane address from CPU
      input  wire [18:35] cpuPC,        // Program counter
      input  wire [ 0:35] cpuHR,        // Instruction register
      input  wire         regsLOAD,     // Load registers
      input  wire         vmaLOAD,      // Load VMA
      input  wire         regTRCMD_WR,  // DCSR trace command write
      input  wire [ 0: 2] regTRCMD,     // DCSR trace command
      input  wire         regBRCMD_WR,  // DCSR breakpoint command write
      input  wire [ 0: 2] regBRCMD,     // DCSR breakpoint command
      output wire [ 0:35] regDCSR,      // DCSR register
      input  wire [ 0:35] regDBAR,      // Breakpoint address register
      input  wire [ 0:35] regDBMR,      // DBAR register
      input  wire         regDITR_RD,   // DITR read
      output wire [ 0:63] regDITR,      // DITR register
      output reg  [ 0:63] regDPCIR,     // DPCIR register
      output wire         debugHALT     // Halt signal to CPU
   );

   //
   // Full/empty flags
   //

   wire trfull;
   wire trempty;

   //
   // Match and mask
   //

   wire match = (cpuADDR & regDBMR) == (regDBAR & regDBMR);

   //
   // Trace Trigger State Machine
   //

   localparam [2:0] regTRCMD_RESET   = 0,
                    regTRCMD_TRIGGER = 1,
                    regTRCMD_ADDRMAT = 2,
                    regTRCMD_STOP    = 3;

   localparam [2:0] trstateIDLE   = 0,
                    trstateARMED  = 1,
                    trstateACTIVE = 2,
                    trstateDONE   = 3;

   reg [2:0] trstate;
   always @(posedge clk or posedge rst)
     begin
        if (rst)
          trstate <= trstateIDLE;
        else
          if ((regTRCMD == regTRCMD_RESET) & regTRCMD_WR)
            trstate <= trstateIDLE;
          else
            case (trstate)
              trstateIDLE:
                if (regTRCMD_WR)
                  case (regTRCMD)
                    regTRCMD_TRIGGER:
                      trstate <= trstateACTIVE;
                    regTRCMD_ADDRMAT:
                      trstate <= trstateARMED;
                  endcase
              trstateARMED:
                if (match)
                  trstate <= trstateACTIVE;
                else if ((regTRCMD == regTRCMD_STOP) & regTRCMD_WR)
                  trstate <= trstateDONE;
              trstateACTIVE:
                if (trfull | ((regTRCMD == regTRCMD_STOP) & regTRCMD_WR))
                  trstate <= trstateDONE;
              trstateDONE:
                trstate <= trstateDONE;
            endcase
     end

   //
   // Breakpoint Trigger State Machine
   //

   localparam [2:0] regBRCMD_DISABLE = 0,
                    regBRCMD_TRIG    = 1,
                    regBRCMD_FULL    = 2,
                    regBRCMD_EITHER  = 3;

   localparam [2:0] brstateIDLE  = 0,
                    brstateARMED = 1,
                    brstateBREAK = 2;

  reg [2:0] brstate;
   always @(posedge clk or posedge rst)
     begin
        if (rst)
          brstate <= trstateIDLE;
        else
          if ((regBRCMD == regBRCMD_DISABLE) & regBRCMD_WR)
            brstate <= brstateIDLE;
          else
            case (brstate)
              brstateIDLE:
                if (regBRCMD_WR)
                  case (regBRCMD)
                    regBRCMD_TRIG,
                    regBRCMD_FULL,
                    regBRCMD_EITHER:
                      brstate <= brstateARMED;
                  endcase
              brstateARMED:
                if (((regBRCMD == regBRCMD_TRIG)   & match ) |
                    ((regBRCMD == regBRCMD_FULL)   & trfull) |
                    ((regBRCMD == regBRCMD_EITHER) & match ) |
                    ((regBRCMD == regBRCMD_EITHER) & trfull))
                  brstate <= brstateBREAK;
              brstateBREAK:
                brstate <= brstateIDLE;
            endcase
     end

   //
   // Instruction Trace Buffer (FIFO)
   //

   wire fifo_rd;
   wire fifo_wr;
   wire [ 0:35] fifoHR;
   wire [18:35] fifoPC;

   EDGETRIG #(
      .POSEDGE    (0)
   ) traceRD (
      .clk        (clk),
      .rst        (rst),
      .clken      (1'b1),
      .i          (regDITR_RD),
      .o          (fifo_rd)
   );

   EDGETRIG #(
      .POSEDGE    (1)
   ) traceWR (
      .clk        (clk),
      .rst        (rst),
      .clken      (1'b1),
      .i          (regsLOAD & (trstate == trstateACTIVE)),
      .o          (fifo_wr)
   );

   FIFO #(
      .SIZE       (16*1024),
      .WIDTH      (54)
   ) TRACE_BUFFER (
      .clk        (clk),
      .rst        (rst),
      .clr        (trstate == trstateIDLE),
      .clken      (1'b1),
      .rd         (fifo_rd),
      .wr         (fifo_wr),
      .in         ({cpuPC, cpuHR}),
      .out        ({fifoPC, fifoHR}),
      .full       (trfull),
      .empty      (trempty)
   );

   //
   // Build Control/Status Register
   //

   assign regDCSR = {12'b0, regBRCMD, brstate, 10'b0, regTRCMD, trstate, trfull, trempty};

   //
   // Build Instruction Trace Register
   //

   assign regDITR = {10'b0, fifoPC, fifoHR};

   //
   // DPCIR Register
   //

   always @(posedge clk or posedge rst)
     begin
        if (rst)
          regDPCIR <= 0;
        else
          if (regsLOAD)
            regDPCIR <= {cpuPC, cpuHR};
     end

   //
   // Breakpoint Halt
   //

   assign debugHALT = brstate == brstateBREAK;

   //
   // Simulation Support
   //
   //  This code is used by the simulator to print the program counter on the
   //  console display as the code executes.   A modified PC does not mean that
   //  the instruction was actually executed.  For example, the PC is always
   //  incremented after the instruction is fetched but the PC may be modified
   //  (again) later by a branch instruction.   This code prints the program
   //  counter when the instruction register is loaded.  This occurs once during
   //  the instruction execution.
   //
   //  This module also has some code that attempts to halt the simulation if
   //  the CPU gets stuck.  It does this by watching for VMA changes and PC
   //  changes.
   //
   //  The PC will appear to be stuck for long period of time when doing BLT
   //  operations therefore watching for just PC changes is not sufficient.
   //

`ifndef SYNTHESIS

   //
   // Registers
   //

   reg [18:35] PC;
   reg [14*8:1] test;

   //
   // Remember last time VMA was updated
   //

   time lastVMA;
   always @(posedge clk or posedge rst)
     begin
        if (rst)
          lastVMA = 0;
        else
          if (vmaLOAD)
            lastVMA = $time;
     end

   //
   // Remember last time IR was updated
   //

   time lastIR;
   always @(posedge clk or posedge rst)
     begin
        if (rst)
          lastIR = 0;
        else
          if (regsLOAD)
            lastIR = $time;

          //
          // Whine if the PC but not the VMA gets stuck for 1 ms
          //

          else if ((($time - lastIR) > 1000000) && (($time - lastVMA) < 1000000))
            begin
               lastIR = $time;
               $display("[%11.3f] %15s: PC is %06o (not stuck).", $time/1.0e3, test, PC);
            end

          //
          // Whine if both the PC and the VMA gets stuck for 1 ms
          //

          else if ((($time - lastIR) > 1000000) && (($time - lastVMA) > 1000000))
            begin
               lastIR = $time;
               $display("[%11.3f] %15s: PC is %06o (stuck).", $time/1.0e3, test, PC);
`ifdef STOP_ON_STUCK_PC
               $stop;
`endif
            end
     end

   //
   // Print out Program Counter in the Simulator
   //

   always @(posedge clk or posedge rst)
     begin
        if (rst)
          begin
             PC   = 0;
             test = "";
          end
        else
          if (regsLOAD)
            begin
               PC     = cpuPC;
               lastIR = $time;

               if (PC == 18'o030057)
                 begin
                    $display("Test Completed.");
`ifdef STOP_ON_COMPLETE
                    $stop;
`endif
                 end

                 `ifdef DEBUG_DSKAH
                    `include "debug_dskah.vh"
                 `elsif DEBUG_DSKBA
                    `include "debug_dskba.vh"
                 `elsif DEBUG_DSKCG
                   `include "debug_dskcg.vh"
                 `elsif DEBUG_DSKEA
                    `include "debug_dskea.vh"
                 `elsif DEBUG_DSKEB
                    `include "debug_dskeb.vh"
                 `elsif DEBUG_DSKEC
                    `include "debug_dskec.vh"
                 `elsif DEBUG_DSDZA
                    `include "debug_dsdza.vh"
                 `elsif DEBUG_DSUBA
                    `include "debug_dsuba.vh"
                 `else
                    `include "debug_default.vh"
                 `endif
                 `include "debug_smmon.vh"

                 $display("[%11.3f] %15s: PC is %06o", $time/1.0e3, test, PC);
            end
     end

`endif

endmodule
