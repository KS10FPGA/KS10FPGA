////////////////////////////////////////////////////////////////////
//!
//! KS-10 Processor
//!
//! \brief
//!      Dispatch ROM (DROM)
//!
//! \details
//!
//! \todo
//!
//! \file
//!      drom.v
//!
//! \author
//!      Rob Doyle - doyle (at) cox (dot) net
//!
////////////////////////////////////////////////////////////////////
//
//  Copyright (C) 2009, 2012 Rob Doyle
//
// This source file may be used and distributed without
// restriction provided that this copyright statement is not
// removed from the file and that any derivative work contains
// the original copyright notice and the associated disclaimer.
//
// This source file is free software; you can redistribute it
// and/or modify it under the terms of the GNU Lesser General
// Public License as published by the Free Software Foundation;
// version 2.1 of the License.
//
// This source is distributed in the hope that it will be
// useful, but WITHOUT ANY WARRANTY; without even the implied
// warranty of MERCHANTABILITY or FITNESS FOR A PARTICULAR
// PURPOSE. See the GNU Lesser General Public License for more
// details.
//
// You should have received a copy of the GNU Lesser General
// Public License along with this source; if not, download it
// from http://www.gnu.org/licenses/lgpl.txt
//
////////////////////////////////////////////////////////////////////
//
// Comments are formatted for doxygen
//

`include "drom.vh"

module DROM(clk, clken, dbus, drom);

   parameter  dromWidth = `DROM_WIDTH;

   input      clk;                  	// Clock
   input      clken;                	// Clock Enable
   input      [0:35]          dbus;   	// Data Bus (Instruction Register)
   output reg [0:dromWidth-1] drom;     // Output Data

   //
   // Dispatch ROM (DROM)
   //  DPEA/E98
   //  DPEA/E117
   //  DPEA/E110
   //

   always @(posedge clk)
     begin
        if (clken)
          case (dbus[0:8])
            //                  0000 1112 2233
            //                  0369 2581 4703
            9'o000: drom <= 36'o0000_1556_2100;
            9'o001: drom <= 36'o0001_1740_2100;
            9'o002: drom <= 36'o0002_1740_2100;
            9'o003: drom <= 36'o0003_1740_2100;
            9'o004: drom <= 36'o0002_1741_2100;
            9'o005: drom <= 36'o0005_1740_2100;
            9'o006: drom <= 36'o0006_1740_2100;
            9'o007: drom <= 36'o0007_1740_2100;
            9'o010: drom <= 36'o0001_1742_2100;
            9'o011: drom <= 36'o0004_1742_2100;
            9'o012: drom <= 36'o0001_1743_2100;
            9'o013: drom <= 36'o0000_1743_2100;
            9'o014: drom <= 36'o0001_1744_2100;
            9'o015: drom <= 36'o0000_1744_2100;
            9'o016: drom <= 36'o0002_1744_2100;
            9'o017: drom <= 36'o0003_1744_2100;
            9'o020: drom <= 36'o0000_1746_2100;
            9'o021: drom <= 36'o0000_1747_2100;
            9'o022: drom <= 36'o0000_1750_2100;
            9'o023: drom <= 36'o0000_1751_2100;
            9'o024: drom <= 36'o0001_1751_2100;
            9'o025: drom <= 36'o0002_1751_2100;
            9'o026: drom <= 36'o0004_1751_2100;
            9'o027: drom <= 36'o0010_1751_2100;
            9'o030: drom <= 36'o0000_1557_2100;
            9'o031: drom <= 36'o0001_1557_2100;
            9'o032: drom <= 36'o0002_1557_2100;
            9'o033: drom <= 36'o0003_1557_2100;
            9'o034: drom <= 36'o0004_1557_2100;
            9'o035: drom <= 36'o0005_1557_2100;
            9'o036: drom <= 36'o0006_1557_2100;
            9'o037: drom <= 36'o0007_1557_2100;
            9'o040: drom <= 36'o0000_1556_2100;
            9'o041: drom <= 36'o0000_1556_2100;
            9'o042: drom <= 36'o0000_1556_2100;
            9'o043: drom <= 36'o0000_1556_2100;
            9'o044: drom <= 36'o0000_1556_2100;
            9'o045: drom <= 36'o0000_1556_2100;
            9'o046: drom <= 36'o0000_1556_2100;
            9'o047: drom <= 36'o0000_1556_2100;
            9'o050: drom <= 36'o0000_1556_2100;
            9'o051: drom <= 36'o0000_1556_2100;
            9'o052: drom <= 36'o0000_1556_2100;
            9'o053: drom <= 36'o0000_1556_2100;
            9'o054: drom <= 36'o0000_1556_2100;
            9'o055: drom <= 36'o0000_1556_2100;
            9'o056: drom <= 36'o0000_1556_2100;
            9'o057: drom <= 36'o0000_1556_2100;
            9'o060: drom <= 36'o0000_1556_2100;
            9'o061: drom <= 36'o0000_1556_2100;
            9'o062: drom <= 36'o0000_1556_2100;
            9'o063: drom <= 36'o0000_1556_2100;
            9'o064: drom <= 36'o0000_1556_2100;
            9'o065: drom <= 36'o0000_1556_2100;
            9'o066: drom <= 36'o0000_1556_2100;
            9'o067: drom <= 36'o0000_1556_2100;
            9'o070: drom <= 36'o0000_1556_2100;
            9'o071: drom <= 36'o0000_1556_2100;
            9'o072: drom <= 36'o0000_1556_2100;
            9'o073: drom <= 36'o0000_1556_2100;
            9'o074: drom <= 36'o0000_1556_2100;
            9'o075: drom <= 36'o0000_1556_2100;
            9'o076: drom <= 36'o0000_1556_2100;
            9'o077: drom <= 36'o0000_1556_2100;
            9'o100: drom <= 36'o0000_1556_2100;
            9'o101: drom <= 36'o0000_1661_2100;
            9'o102: drom <= 36'o0000_1662_2100;
            9'o103: drom <= 36'o0000_1663_2100;
            9'o104: drom <= 36'o0000_1664_2100;
            9'o105: drom <= 36'o0000_1551_3000;
            9'o106: drom <= 36'o0000_1666_2100;
            9'o107: drom <= 36'o0000_1667_2100;
            9'o110: drom <= 36'o1100_1637_1100;
            9'o111: drom <= 36'o1100_1635_1100;
            9'o112: drom <= 36'o1105_1631_1100;
            9'o113: drom <= 36'o1105_1636_1100;
            9'o114: drom <= 36'o0205_1457_1100;
            9'o115: drom <= 36'o0205_1615_1100;
            9'o116: drom <= 36'o0205_1566_1100;
            9'o117: drom <= 36'o0205_1627_1100;
            9'o120: drom <= 36'o0205_1505_1100;
            9'o121: drom <= 36'o0215_1434_1100;
            9'o122: drom <= 36'o0701_1626_1100;
            9'o123: drom <= 36'o0000_1467_3100;
            9'o124: drom <= 36'o0300_1567_0100;
            9'o125: drom <= 36'o0100_1565_0500;
            9'o126: drom <= 36'o0711_1626_1100;
            9'o127: drom <= 36'o0011_1616_1100;
            9'o130: drom <= 36'o0000_1660_2100;
            9'o131: drom <= 36'o0001_1660_2100;
            9'o132: drom <= 36'o0001_1621_2100;
            9'o133: drom <= 36'o0015_1610_1100;
            9'o134: drom <= 36'o0000_1620_1500;
            9'o135: drom <= 36'o0000_1624_1100;
            9'o136: drom <= 36'o0000_1630_1500;
            9'o137: drom <= 36'o0000_1634_1100;
            9'o140: drom <= 36'o0701_1577_1100;
            9'o141: drom <= 36'o0002_1660_2100;
            9'o142: drom <= 36'o0702_1577_1700;
            9'o143: drom <= 36'o0703_1577_1700;
            9'o144: drom <= 36'o0711_1577_1100;
            9'o145: drom <= 36'o0611_1577_0100;
            9'o146: drom <= 36'o0712_1577_1700;
            9'o147: drom <= 36'o0713_1577_1700;
            9'o150: drom <= 36'o0701_1576_1100;
            9'o151: drom <= 36'o0003_1660_2100;
            9'o152: drom <= 36'o0702_1576_1700;
            9'o153: drom <= 36'o0703_1576_1700;
            9'o154: drom <= 36'o0711_1576_1100;
            9'o155: drom <= 36'o0611_1576_0100;
            9'o156: drom <= 36'o0712_1576_1700;
            9'o157: drom <= 36'o0713_1576_1700;
            9'o160: drom <= 36'o0701_1570_1100;
            9'o161: drom <= 36'o0004_1660_2100;
            9'o162: drom <= 36'o0702_1570_1700;
            9'o163: drom <= 36'o0703_1570_1700;
            9'o164: drom <= 36'o0711_1570_1100;
            9'o165: drom <= 36'o0611_1570_0100;
            9'o166: drom <= 36'o0712_1570_1700;
            9'o167: drom <= 36'o0713_1570_1700;
            9'o170: drom <= 36'o0701_1574_1100;
            9'o171: drom <= 36'o0005_1660_2100;
            9'o172: drom <= 36'o0702_1574_1700;
            9'o173: drom <= 36'o0703_1574_1700;
            9'o174: drom <= 36'o0711_1574_1100;
            9'o175: drom <= 36'o0611_1574_0100;
            9'o176: drom <= 36'o0712_1574_1700;
            9'o177: drom <= 36'o0713_1574_1700;
            9'o200: drom <= 36'o1015_1515_1100;
            9'o201: drom <= 36'o0015_1515_3000;
            9'o202: drom <= 36'o0116_1404_0700;
            9'o203: drom <= 36'o0004_1504_1700;
            9'o204: drom <= 36'o1015_1402_1100;
            9'o205: drom <= 36'o0015_1402_3000;
            9'o206: drom <= 36'o0116_1402_0700;
            9'o207: drom <= 36'o0004_1402_1700;
            9'o210: drom <= 36'o1015_1405_1100;
            9'o211: drom <= 36'o0015_1405_3000;
            9'o212: drom <= 36'o0116_1405_0700;
            9'o213: drom <= 36'o0004_1405_1700;
            9'o214: drom <= 36'o1015_1403_1100;
            9'o215: drom <= 36'o0015_1515_3000;
            9'o216: drom <= 36'o0116_1403_0700;
            9'o217: drom <= 36'o0004_1403_1700;
            9'o220: drom <= 36'o1015_1641_1100;
            9'o221: drom <= 36'o0015_1641_3000;
            9'o222: drom <= 36'o0016_1641_1700;
            9'o223: drom <= 36'o0017_1641_1700;
            9'o224: drom <= 36'o1005_1571_1100;
            9'o225: drom <= 36'o0005_1571_3000;
            9'o226: drom <= 36'o0016_1571_1700;
            9'o227: drom <= 36'o0006_1571_1700;
            9'o230: drom <= 36'o1005_1600_1100;
            9'o231: drom <= 36'o0005_1600_3000;
            9'o232: drom <= 36'o0016_1600_1700;
            9'o233: drom <= 36'o0006_1600_1700;
            9'o234: drom <= 36'o1005_1601_1100;
            9'o235: drom <= 36'o0005_1601_3000;
            9'o236: drom <= 36'o0016_1601_1700;
            9'o237: drom <= 36'o0006_1601_1700;
            9'o240: drom <= 36'o0400_1622_1000;
            9'o241: drom <= 36'o0400_1632_1000;
            9'o242: drom <= 36'o0400_1612_1000;
            9'o243: drom <= 36'o0000_1462_2100;
            9'o244: drom <= 36'o0000_1466_3000;
            9'o245: drom <= 36'o0500_1470_1000;
            9'o246: drom <= 36'o0500_1464_1000;
            9'o247: drom <= 36'o0000_1665_2100;
            9'o250: drom <= 36'o0015_1406_1500;
            9'o251: drom <= 36'o0000_1640_2100;
            9'o252: drom <= 36'o0005_1547_2100;
            9'o253: drom <= 36'o0001_1547_2100;
            9'o254: drom <= 36'o0000_1520_6000;
            9'o255: drom <= 36'o0000_1540_2100;
            9'o256: drom <= 36'o0000_1541_1100;
            9'o257: drom <= 36'o1215_1553_0100;
            9'o260: drom <= 36'o0000_1544_2100;
            9'o261: drom <= 36'o0002_1543_3100;
            9'o262: drom <= 36'o0002_1545_2100;
            9'o263: drom <= 36'o0000_1546_2100;
            9'o264: drom <= 36'o0000_1552_2100;
            9'o265: drom <= 36'o0000_1550_2100;
            9'o266: drom <= 36'o0000_1554_2100;
            9'o267: drom <= 36'o0000_1555_2100;
            9'o270: drom <= 36'o1015_1560_1100;
            9'o271: drom <= 36'o0015_1560_3000;
            9'o272: drom <= 36'o0016_1560_1700;
            9'o273: drom <= 36'o0017_1560_1700;
            9'o274: drom <= 36'o1015_1561_1100;
            9'o275: drom <= 36'o0015_1561_3000;
            9'o276: drom <= 36'o0016_1561_1700;
            9'o277: drom <= 36'o0017_1561_1700;
            9'o300: drom <= 36'o0000_1400_2100;
            9'o301: drom <= 36'o0001_1476_2100;
            9'o302: drom <= 36'o0002_1476_2100;
            9'o303: drom <= 36'o0003_1476_2100;
            9'o304: drom <= 36'o0004_1476_2100;
            9'o305: drom <= 36'o0005_1476_2100;
            9'o306: drom <= 36'o0006_1476_2100;
            9'o307: drom <= 36'o0007_1476_2100;
            9'o310: drom <= 36'o0000_1476_1100;
            9'o311: drom <= 36'o0001_1476_1100;
            9'o312: drom <= 36'o0002_1476_1100;
            9'o313: drom <= 36'o0003_1476_1100;
            9'o314: drom <= 36'o0004_1476_1100;
            9'o315: drom <= 36'o0005_1476_1100;
            9'o316: drom <= 36'o0006_1476_1100;
            9'o317: drom <= 36'o0007_1476_1100;
            9'o320: drom <= 36'o0000_1400_2100;
            9'o321: drom <= 36'o0001_1440_2100;
            9'o322: drom <= 36'o0002_1440_2100;
            9'o323: drom <= 36'o0003_1440_2100;
            9'o324: drom <= 36'o0004_1520_2100;
            9'o325: drom <= 36'o0005_1440_2100;
            9'o326: drom <= 36'o0006_1440_2100;
            9'o327: drom <= 36'o0007_1440_2100;
            9'o330: drom <= 36'o0000_1477_1100;
            9'o331: drom <= 36'o0001_1477_1100;
            9'o332: drom <= 36'o0002_1477_1100;
            9'o333: drom <= 36'o0003_1477_1100;
            9'o334: drom <= 36'o0004_1477_1100;
            9'o335: drom <= 36'o0005_1477_1100;
            9'o336: drom <= 36'o0006_1477_1100;
            9'o337: drom <= 36'o0007_1477_1100;
            9'o340: drom <= 36'o0000_1611_3000;
            9'o341: drom <= 36'o0001_1611_2100;
            9'o342: drom <= 36'o0002_1611_2100;
            9'o343: drom <= 36'o0003_1611_2100;
            9'o344: drom <= 36'o0004_1611_2100;
            9'o345: drom <= 36'o0005_1611_2100;
            9'o346: drom <= 36'o0006_1611_2100;
            9'o347: drom <= 36'o0007_1611_2100;
            9'o350: drom <= 36'o0000_1431_1500;
            9'o351: drom <= 36'o0001_1431_1500;
            9'o352: drom <= 36'o0002_1431_1500;
            9'o353: drom <= 36'o0003_1431_1500;
            9'o354: drom <= 36'o0004_1431_1500;
            9'o355: drom <= 36'o0005_1431_1500;
            9'o356: drom <= 36'o0006_1431_1500;
            9'o357: drom <= 36'o0007_1431_1500;
            9'o360: drom <= 36'o0000_1542_3000;
            9'o361: drom <= 36'o0001_1542_2100;
            9'o362: drom <= 36'o0002_1542_2100;
            9'o363: drom <= 36'o0003_1542_2100;
            9'o364: drom <= 36'o0004_1542_2100;
            9'o365: drom <= 36'o0005_1542_2100;
            9'o366: drom <= 36'o0006_1542_2100;
            9'o367: drom <= 36'o0007_1542_2100;
            9'o370: drom <= 36'o0000_1437_1500;
            9'o371: drom <= 36'o0001_1437_1500;
            9'o372: drom <= 36'o0002_1437_1500;
            9'o373: drom <= 36'o0003_1437_1500;
            9'o374: drom <= 36'o0004_1437_1500;
            9'o375: drom <= 36'o0005_1437_1500;
            9'o376: drom <= 36'o0006_1437_1500;
            9'o377: drom <= 36'o0007_1437_1500;
            9'o400: drom <= 36'o0015_1441_3000;
            9'o401: drom <= 36'o0015_1441_3000;
            9'o402: drom <= 36'o0016_1441_2700;
            9'o403: drom <= 36'o0017_1441_2700;
            9'o404: drom <= 36'o1015_1442_1100;
            9'o405: drom <= 36'o0015_1442_3000;
            9'o406: drom <= 36'o0016_1442_1700;
            9'o407: drom <= 36'o0017_1442_1700;
            9'o410: drom <= 36'o1015_1443_1100;
            9'o411: drom <= 36'o0015_1443_3000;
            9'o412: drom <= 36'o0016_1443_1700;
            9'o413: drom <= 36'o0017_1443_1700;
            9'o414: drom <= 36'o1015_1404_1100;
            9'o415: drom <= 36'o0015_1404_3000;
            9'o416: drom <= 36'o0016_1404_1700;
            9'o417: drom <= 36'o0017_1404_1700;
            9'o420: drom <= 36'o1015_1444_1100;
            9'o421: drom <= 36'o0015_1444_3000;
            9'o422: drom <= 36'o0016_1444_1700;
            9'o423: drom <= 36'o0017_1444_1700;
            9'o424: drom <= 36'o0000_1400_1100;
            9'o425: drom <= 36'o0000_1400_2100;
            9'o426: drom <= 36'o0116_1404_0700;
            9'o427: drom <= 36'o0116_1404_0700;
            9'o430: drom <= 36'o1015_1445_1100;
            9'o431: drom <= 36'o0015_1445_3000;
            9'o432: drom <= 36'o0016_1445_1700;
            9'o433: drom <= 36'o0017_1445_1700;
            9'o434: drom <= 36'o1015_1446_1100;
            9'o435: drom <= 36'o0015_1446_3000;
            9'o436: drom <= 36'o0016_1446_1700;
            9'o437: drom <= 36'o0017_1446_1700;
            9'o440: drom <= 36'o1015_1447_1100;
            9'o441: drom <= 36'o0015_1447_3000;
            9'o442: drom <= 36'o0016_1447_1700;
            9'o443: drom <= 36'o0017_1447_1700;
            9'o444: drom <= 36'o1015_1450_1100;
            9'o445: drom <= 36'o0015_1450_3000;
            9'o446: drom <= 36'o0016_1450_1700;
            9'o447: drom <= 36'o0017_1450_1700;
            9'o450: drom <= 36'o0015_1451_3000;
            9'o451: drom <= 36'o0015_1451_3000;
            9'o452: drom <= 36'o0016_1451_2700;
            9'o453: drom <= 36'o0017_1451_2700;
            9'o454: drom <= 36'o1015_1452_1100;
            9'o455: drom <= 36'o0015_1452_3000;
            9'o456: drom <= 36'o0016_1452_1700;
            9'o457: drom <= 36'o0017_1452_1700;
            9'o460: drom <= 36'o1015_1453_1100;
            9'o461: drom <= 36'o0015_1453_3000;
            9'o462: drom <= 36'o0016_1453_1700;
            9'o463: drom <= 36'o0017_1453_1700;
            9'o464: drom <= 36'o1015_1454_1100;
            9'o465: drom <= 36'o0015_1454_3000;
            9'o466: drom <= 36'o0016_1454_1700;
            9'o467: drom <= 36'o0017_1454_1700;
            9'o470: drom <= 36'o1015_1455_1100;
            9'o471: drom <= 36'o0015_1455_3000;
            9'o472: drom <= 36'o0016_1455_1700;
            9'o473: drom <= 36'o0017_1455_1700;
            9'o474: drom <= 36'o0015_1456_3000;
            9'o475: drom <= 36'o0015_1456_3000;
            9'o476: drom <= 36'o0016_1456_2700;
            9'o477: drom <= 36'o0017_1456_2700;
            9'o500: drom <= 36'o1015_1410_1100;
            9'o501: drom <= 36'o0015_1410_3000;
            9'o502: drom <= 36'o0016_1407_1700;
            9'o503: drom <= 36'o0004_1404_1700;
            9'o504: drom <= 36'o1015_1411_1100;
            9'o505: drom <= 36'o0015_1411_3000;
            9'o506: drom <= 36'o0016_1413_1700;
            9'o507: drom <= 36'o0004_1414_1700;
            9'o510: drom <= 36'o1015_1432_1100;
            9'o511: drom <= 36'o0015_1432_3000;
            9'o512: drom <= 36'o0116_1432_0700;
            9'o513: drom <= 36'o0004_1432_1700;
            9'o514: drom <= 36'o1015_1424_1100;
            9'o515: drom <= 36'o0015_1424_3000;
            9'o516: drom <= 36'o0116_1424_0700;
            9'o517: drom <= 36'o0004_1424_1700;
            9'o520: drom <= 36'o1015_1433_1100;
            9'o521: drom <= 36'o0015_1433_3000;
            9'o522: drom <= 36'o0116_1433_0700;
            9'o523: drom <= 36'o0004_1433_1700;
            9'o524: drom <= 36'o1015_1425_1100;
            9'o525: drom <= 36'o0015_1425_3000;
            9'o526: drom <= 36'o0116_1425_0700;
            9'o527: drom <= 36'o0004_1425_1700;
            9'o530: drom <= 36'o1015_1430_1100;
            9'o531: drom <= 36'o0015_1430_3000;
            9'o532: drom <= 36'o0116_1430_0700;
            9'o533: drom <= 36'o0004_1430_1700;
            9'o534: drom <= 36'o1015_1422_1100;
            9'o535: drom <= 36'o0015_1422_3000;
            9'o536: drom <= 36'o0116_1422_0700;
            9'o537: drom <= 36'o0004_1422_1700;
            9'o540: drom <= 36'o1015_1407_1100;
            9'o541: drom <= 36'o0015_1407_3000;
            9'o542: drom <= 36'o0016_1410_1700;
            9'o543: drom <= 36'o0004_1404_1700;
            9'o544: drom <= 36'o1015_1412_1100;
            9'o545: drom <= 36'o0015_1412_3000;
            9'o546: drom <= 36'o0016_1415_1700;
            9'o547: drom <= 36'o0004_1416_1700;
            9'o550: drom <= 36'o1015_1420_1100;
            9'o551: drom <= 36'o0015_1420_3000;
            9'o552: drom <= 36'o0116_1420_0700;
            9'o553: drom <= 36'o0004_1420_1700;
            9'o554: drom <= 36'o1015_1426_1100;
            9'o555: drom <= 36'o0015_1426_3000;
            9'o556: drom <= 36'o0116_1426_0700;
            9'o557: drom <= 36'o0004_1426_1700;
            9'o560: drom <= 36'o1015_1421_1100;
            9'o561: drom <= 36'o0015_1421_3000;
            9'o562: drom <= 36'o0116_1421_0700;
            9'o563: drom <= 36'o0004_1421_1700;
            9'o564: drom <= 36'o1015_1427_1100;
            9'o565: drom <= 36'o0015_1427_3000;
            9'o566: drom <= 36'o0116_1427_0700;
            9'o567: drom <= 36'o0004_1427_1700;
            9'o570: drom <= 36'o1015_1417_1100;
            9'o571: drom <= 36'o0015_1417_3000;
            9'o572: drom <= 36'o0116_1417_0700;
            9'o573: drom <= 36'o0004_1417_1700;
            9'o574: drom <= 36'o1015_1423_1100;
            9'o575: drom <= 36'o0015_1423_3000;
            9'o576: drom <= 36'o0116_1423_0700;
            9'o577: drom <= 36'o0004_1423_1700;
            9'o600: drom <= 36'o0000_1400_2100;
            9'o601: drom <= 36'o0000_1400_2100;
            9'o602: drom <= 36'o0000_1475_2100;
            9'o603: drom <= 36'o0000_1474_2100;
            9'o604: drom <= 36'o0000_1473_2100;
            9'o605: drom <= 36'o0000_1472_2100;
            9'o606: drom <= 36'o0004_1475_2100;
            9'o607: drom <= 36'o0004_1474_2100;
            9'o610: drom <= 36'o0000_1400_2100;
            9'o611: drom <= 36'o0000_1400_2100;
            9'o612: drom <= 36'o0000_1475_1100;
            9'o613: drom <= 36'o0000_1474_1100;
            9'o614: drom <= 36'o0000_1473_1100;
            9'o615: drom <= 36'o0000_1472_1100;
            9'o616: drom <= 36'o0004_1475_1100;
            9'o617: drom <= 36'o0004_1474_1100;
            9'o620: drom <= 36'o0005_1473_2100;
            9'o621: drom <= 36'o0005_1472_2100;
            9'o622: drom <= 36'o0001_1475_2100;
            9'o623: drom <= 36'o0001_1474_2100;
            9'o624: drom <= 36'o0001_1473_2100;
            9'o625: drom <= 36'o0001_1472_2100;
            9'o626: drom <= 36'o0005_1475_2100;
            9'o627: drom <= 36'o0005_1474_2100;
            9'o630: drom <= 36'o0005_1473_1100;
            9'o631: drom <= 36'o0005_1472_1100;
            9'o632: drom <= 36'o0001_1475_1100;
            9'o633: drom <= 36'o0001_1474_1100;
            9'o634: drom <= 36'o0001_1473_1100;
            9'o635: drom <= 36'o0001_1472_1100;
            9'o636: drom <= 36'o0005_1475_1100;
            9'o637: drom <= 36'o0005_1474_1100;
            9'o640: drom <= 36'o0006_1473_2100;
            9'o641: drom <= 36'o0006_1472_2100;
            9'o642: drom <= 36'o0002_1475_2100;
            9'o643: drom <= 36'o0002_1474_2100;
            9'o644: drom <= 36'o0002_1473_2100;
            9'o645: drom <= 36'o0002_1472_2100;
            9'o646: drom <= 36'o0006_1475_2100;
            9'o647: drom <= 36'o0006_1474_2100;
            9'o650: drom <= 36'o0006_1473_1100;
            9'o651: drom <= 36'o0006_1472_1100;
            9'o652: drom <= 36'o0002_1475_1100;
            9'o653: drom <= 36'o0002_1474_1100;
            9'o654: drom <= 36'o0002_1473_1100;
            9'o655: drom <= 36'o0002_1472_1100;
            9'o656: drom <= 36'o0006_1475_1100;
            9'o657: drom <= 36'o0006_1474_1100;
            9'o660: drom <= 36'o0007_1473_2100;
            9'o661: drom <= 36'o0007_1472_2100;
            9'o662: drom <= 36'o0003_1475_2100;
            9'o663: drom <= 36'o0003_1474_2100;
            9'o664: drom <= 36'o0003_1473_2100;
            9'o665: drom <= 36'o0003_1472_2100;
            9'o666: drom <= 36'o0007_1475_2100;
            9'o667: drom <= 36'o0007_1474_2100;
            9'o670: drom <= 36'o0007_1473_1100;
            9'o671: drom <= 36'o0007_1472_1100;
            9'o672: drom <= 36'o0003_1475_1100;
            9'o673: drom <= 36'o0003_1474_1100;
            9'o674: drom <= 36'o0003_1473_1100;
            9'o675: drom <= 36'o0003_1472_1100;
            9'o676: drom <= 36'o0007_1475_1100;
            9'o677: drom <= 36'o0007_1474_1100;
            9'o700: drom <= 36'o1200_1700_4100;
            9'o701: drom <= 36'o1200_1720_4100;
            9'o702: drom <= 36'o1216_1760_4700;
            9'o703: drom <= 36'o0003_1650_2100;
            9'o704: drom <= 36'o1200_1754_0100;
            9'o705: drom <= 36'o1200_1755_0100;
            9'o706: drom <= 36'o0006_1650_2100;
            9'o707: drom <= 36'o0007_1650_2100;
            9'o710: drom <= 36'o1210_1614_0100;
            9'o711: drom <= 36'o1214_1614_0100;
            9'o712: drom <= 36'o1210_1460_0100;
            9'o713: drom <= 36'o1210_1461_0100;
            9'o714: drom <= 36'o1210_1644_0100;
            9'o715: drom <= 36'o1214_1644_0100;
            9'o716: drom <= 36'o0006_1651_2100;
            9'o717: drom <= 36'o0007_1651_2100;
            9'o720: drom <= 36'o1200_1614_0100;
            9'o721: drom <= 36'o1204_1614_0100;
            9'o722: drom <= 36'o1200_1460_0100;
            9'o723: drom <= 36'o1200_1461_0100;
            9'o724: drom <= 36'o1200_1644_0100;
            9'o725: drom <= 36'o1204_1644_0100;
            9'o726: drom <= 36'o0006_1652_2100;
            9'o727: drom <= 36'o0007_1652_2100;
            9'o730: drom <= 36'o0000_1653_2100;
            9'o731: drom <= 36'o0001_1653_2100;
            9'o732: drom <= 36'o0002_1653_2100;
            9'o733: drom <= 36'o0003_1653_2100;
            9'o734: drom <= 36'o0004_1653_2100;
            9'o735: drom <= 36'o0005_1653_2100;
            9'o736: drom <= 36'o0006_1653_2100;
            9'o737: drom <= 36'o0007_1653_2100;
            9'o740: drom <= 36'o0000_1654_2100;
            9'o741: drom <= 36'o0001_1654_2100;
            9'o742: drom <= 36'o0002_1654_2100;
            9'o743: drom <= 36'o0003_1654_2100;
            9'o744: drom <= 36'o0004_1654_2100;
            9'o745: drom <= 36'o0005_1654_2100;
            9'o746: drom <= 36'o0006_1654_2100;
            9'o747: drom <= 36'o0007_1654_2100;
            9'o750: drom <= 36'o0000_1655_2100;
            9'o751: drom <= 36'o0001_1655_2100;
            9'o752: drom <= 36'o0002_1655_2100;
            9'o753: drom <= 36'o0003_1655_2100;
            9'o754: drom <= 36'o0004_1655_2100;
            9'o755: drom <= 36'o0005_1655_2100;
            9'o756: drom <= 36'o0006_1655_2100;
            9'o757: drom <= 36'o0007_1655_2100;
            9'o760: drom <= 36'o0000_1656_2100;
            9'o761: drom <= 36'o0001_1656_2100;
            9'o762: drom <= 36'o0002_1656_2100;
            9'o763: drom <= 36'o0003_1656_2100;
            9'o764: drom <= 36'o0004_1656_2100;
            9'o765: drom <= 36'o0005_1656_2100;
            9'o766: drom <= 36'o0006_1656_2100;
            9'o767: drom <= 36'o0007_1656_2100;
            9'o770: drom <= 36'o0000_1657_2100;
            9'o771: drom <= 36'o0001_1657_2100;
            9'o772: drom <= 36'o0002_1657_2100;
            9'o773: drom <= 36'o0003_1657_2100;
            9'o774: drom <= 36'o0004_1657_2100;
            9'o775: drom <= 36'o0005_1657_2100;
            9'o776: drom <= 36'o0006_1657_2100;
            9'o777: drom <= 36'o0007_1657_2100;
          endcase
     end

endmodule
