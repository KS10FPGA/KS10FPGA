////////////////////////////////////////////////////////////////////////////////
//
// KS-10 Processor
//
// Brief
//   LP20 Page Count Register (PCTR)
//
// Details
//   The module implements the LP20 PCTR Register.
//
// File
//   lppctr.v
//
// Author
//   Rob Doyle - doyle (at) cox (dot) net
//
////////////////////////////////////////////////////////////////////////////////
//
// Copyright (C) 2012-2016 Rob Doyle
//
// This source file may be used and distributed without restriction provided
// that this copyright statement is not removed from the file and that any
// derivative work contains the original copyright notice and the associated
// disclaimer.
//
// This source file is free software; you can redistribute it and/or modify it
// under the terms of the GNU Lesser General Public License as published by the
// Free Software Foundation; version 2.1 of the License.
//
// This source is distributed in the hope that it will be useful, but WITHOUT
// ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
// FITNESS FOR A PARTICULAR PURPOSE. See the GNU Lesser General Public License
// for more details.
//
// You should have received a copy of the GNU Lesser General Public License
// along with this source; if not, download it from
// http://www.gnu.org/licenses/lgpl.txt
//
////////////////////////////////////////////////////////////////////////////////

`default_nettype none
`timescale 1ns/1ps

`include "lppctr.vh"

module LPPCTR (
      input  wire         clk,                  // Clock
      input  wire         rst,                  // Reset
      input  wire [35: 0] lpDATAI,              // Bus data in
      input  wire         pctrWRITE,            // Write to PCTR
      input  wire         lpINIT,               // Initialize
      input  wire         lpDECPCTR,            // Decrement PCTR
      output wire         lpPCZ,                // Page counter is zero
      output wire [15: 0] regPCTR               // PCTR output
   );

   //
   // Page count register
   //
   // Trace
   //  M8597/LPD4/E22
   //  M8597/LPD4/E30
   //  M8597/LPD4/E38
   //

   reg [11:0] count;
   always @(posedge clk or posedge rst)
     begin
        if (rst)
          count <= 0;
        else
          begin
             if (lpINIT)
               count <= 0;
             else if (pctrWRITE)
               count <= `lpPCTR_DAT(lpDATAI);
             else if (lpDECPCTR)
               count <= count - 1'b1;
          end
     end

   //
   // Build PCTR Register
   //

   assign regPCTR = {4'b0, count};

   //
   // Page counter is zero
   //
   // Trace
   //  M8597/LPD4/E38
   //

   assign lpPCZ = (count == 0);

endmodule
