////////////////////////////////////////////////////////////////////
//!
//! KS-10 Processor
//!
//! \brief
//!      Microcontroller Control ROM 
//!
//! \details
//!
//! \todo
//!
//! \file
//!      crom.v
//!
//! \author
//!      Rob Doyle - doyle (at) cox (dot) net
//!
////////////////////////////////////////////////////////////////////
//
//  Copyright (C) 2009, 2012 Rob Doyle
//
// This source file may be used and distributed without
// restriction provided that this copyright statement is not
// removed from the file and that any derivative work contains
// the original copyright notice and the associated disclaimer.
//
// This source file is free software; you can redistribute it
// and/or modify it under the terms of the GNU Lesser General
// Public License as published by the Free Software Foundation;
// version 2.1 of the License.
//
// This source is distributed in the hope that it will be
// useful, but WITHOUT ANY WARRANTY; without even the implied
// warranty of MERCHANTABILITY or FITNESS FOR A PARTICULAR
// PURPOSE. See the GNU Lesser General Public License for more
// details.
//
// You should have received a copy of the GNU Lesser General
// Public License along with this source; if not, download it
// from http://www.gnu.org/licenses/lgpl.txt
//
////////////////////////////////////////////////////////////////////
//
// Comments are formatted for doxygen
//

`include "crom.vh"

module CROM(clk, clken, addr, crom);

   parameter  cromWidth = `CROM_WIDTH;
   
   input      clk;                  	// Clock
   input      clken;                	// Clock Enable
   input      [0:11] addr;          	// Address
   output reg [0:cromWidth-1] crom; 	// Output Data 

   //
   // CROM
   //   Note ROM MSB is ignored.
   //
   
   always @(posedge clk)
     begin
        if (clken)
	  case(addr[1:11])
            //                                                               11
            //                     0000 1112 2233 3344 4555 6666 7778 8899 9900
            //                     0369 2581 4703 6925 8147 0369 2581 4703 6925 
            12'o0000: crom <= 108'o0002_3771_0012_4374_4007_0700_0000_0037_7777;
            12'o0001: crom <= 108'o3676_3333_0004_7174_4007_0700_0410_0000_0212;
            12'o0002: crom <= 108'o0013_3445_1212_4174_4007_0700_0000_0000_0000;
            12'o0003: crom <= 108'o0100_4751_1203_4374_4007_0700_0000_0037_6000;
            12'o0004: crom <= 108'o2476_4443_0000_4174_4107_0640_0000_0000_0062;
            12'o0005: crom <= 108'o0004_4443_0000_4174_4007_0660_0000_0000_0000;
            12'o0006: crom <= 108'o3412_4443_0000_4174_4007_0700_0010_0000_0000;
            12'o0007: crom <= 108'o3423_4443_0000_4174_4007_0700_0000_0000_0000;
            12'o0010: crom <= 108'o0560_3771_0004_1276_6007_0701_0010_0000_1444;
            12'o0011: crom <= 108'o0024_3771_0004_7274_4007_0701_0000_0000_0227;
            12'o0012: crom <= 108'o0324_3333_0005_6174_4007_0700_0400_0000_0000;
            12'o0013: crom <= 108'o0053_3551_1212_4374_4007_0700_0000_0000_0001;
            12'o0014: crom <= 108'o1400_3333_0005_4174_4007_0571_0000_0000_0000;
            12'o0015: crom <= 108'o1116_7441_0303_4174_4007_0700_0000_0000_0000;
            12'o0016: crom <= 108'o1123_6551_0303_0274_4007_0700_0000_0000_0000;
            12'o0017: crom <= 108'o1123_3551_0303_0274_4007_0700_0000_0000_0000;
            12'o0020: crom <= 108'o2746_4221_0002_4174_0007_0700_0010_0000_0000;
            12'o0021: crom <= 108'o3000_3446_0606_4174_4007_0700_0010_0000_0000;
            12'o0022: crom <= 108'o3541_3333_0002_4175_5007_0701_0210_0000_0002;
            12'o0023: crom <= 108'o3667_0111_0704_4170_4007_0700_0210_0023_1016;
            12'o0024: crom <= 108'o3700_4223_0000_4364_4277_0700_0210_0000_0010;
            12'o0025: crom <= 108'o1176_3333_0004_4174_4007_0621_0000_0000_0000;
            12'o0026: crom <= 108'o2475_4443_0000_4174_4107_0700_0000_0000_0074;
            12'o0027: crom <= 108'o2740_4751_1205_4374_4007_0700_0000_0000_0430;
            12'o0030: crom <= 108'o0002_3773_0000_2274_4464_1700_0000_0001_0004;
            12'o0031: crom <= 108'o3000_3446_0606_4174_4007_0700_0010_0000_0000;
            12'o0032: crom <= 108'o0002_3333_0002_4174_4464_1700_0000_0001_0004;
            12'o0033: crom <= 108'o3060_4443_0000_4174_4007_0700_0010_0000_0000;
            12'o0034: crom <= 108'o2556_0551_0202_2270_4007_0700_0200_0004_0012;
            12'o0035: crom <= 108'o2760_3445_0403_4174_4007_0700_0000_0000_0000;
            12'o0036: crom <= 108'o2556_3443_0200_4174_4007_0700_0200_0004_0112;
            12'o0037: crom <= 108'o0555_4443_0000_4174_4467_0700_0000_0051_1000;
            12'o0040: crom <= 108'o0000_3771_0003_4365_5001_2700_0200_0000_0002;
            12'o0041: crom <= 108'o0000_3771_0003_0276_6001_2700_0000_0000_0000;
            12'o0042: crom <= 108'o0401_3771_0003_4365_5007_0700_0200_0000_0002;
            12'o0043: crom <= 108'o0415_3771_0003_0276_6007_0700_0000_0000_0000;
            12'o0044: crom <= 108'o0000_3333_0003_4174_4001_2530_3000_0041_5777;
            12'o0045: crom <= 108'o0416_3772_0000_1275_5007_0701_0000_0000_1441;
            12'o0046: crom <= 108'o0372_3770_0303_4344_4007_0700_0000_0000_0000;
            12'o0047: crom <= 108'o0372_3771_0003_4365_5007_0700_0200_0000_0002;
            12'o0050: crom <= 108'o0000_3770_0103_4365_5001_2700_0200_0014_0012;
            12'o0051: crom <= 108'o0402_3771_0005_4365_5177_0521_3000_0041_2000;
            12'o0052: crom <= 108'o0404_4443_0000_4174_4007_0040_0000_0000_0000;
            12'o0053: crom <= 108'o0061_3447_1200_4174_4007_0700_0000_0000_0000;
            12'o0054: crom <= 108'o1232_4552_0000_1275_5007_0701_0000_0000_1441;
            12'o0055: crom <= 108'o3060_6551_1717_4374_4007_0700_0010_0000_0007;
            12'o0056: crom <= 108'o3027_0001_1616_4174_4007_0700_0000_0000_0000;
            12'o0057: crom <= 108'o3025_2225_0016_4174_4007_0700_4000_0000_0000;
            12'o0060: crom <= 108'o3667_3443_0300_4174_4007_0700_0210_0003_0012;
            12'o0061: crom <= 108'o0071_3771_0015_4374_4007_0700_0000_0000_0001;
            12'o0062: crom <= 108'o3000_3446_0606_4174_4007_0700_0010_0000_0000;
            12'o0063: crom <= 108'o1372_3333_0003_4174_4007_0520_0000_0000_0000;
            12'o0064: crom <= 108'o3670_0111_0703_4170_4007_0700_0210_0003_0012;
            12'o0065: crom <= 108'o2606_0111_0703_4174_4007_0700_0200_0004_0002;
            12'o0066: crom <= 108'o3147_0661_0003_7274_4007_0701_0000_0000_0225;
            12'o0067: crom <= 108'o2440_4571_1205_4374_4007_0700_0000_0024_1220;
            12'o0070: crom <= 108'o3101_0553_0300_2274_4007_0700_0200_0004_0712;
            12'o0071: crom <= 108'o0003_4751_1207_4374_4007_0700_0010_0000_0001;
            12'o0072: crom <= 108'o3101_3443_0300_4174_4007_0700_0200_0004_0712;
            12'o0073: crom <= 108'o1514_0111_0503_4174_4003_7700_0200_0003_0001;
            12'o0074: crom <= 108'o3100_0553_0300_2274_4007_0700_0200_0004_0512;
            12'o0075: crom <= 108'o0054_3447_0303_4174_4007_0700_0000_0000_0000;
            12'o0076: crom <= 108'o3100_3443_0300_4174_4007_0700_0200_0004_0512;
            12'o0077: crom <= 108'o2440_4571_1205_4374_4007_0700_0000_0024_1200;
            12'o0100: crom <= 108'o0106_3333_0003_7174_4007_0700_0400_0000_0227;
            12'o0101: crom <= 108'o3474_4751_1203_4374_4367_0700_0000_0000_0423;
            12'o0102: crom <= 108'o3474_4751_1203_4374_4367_0700_0000_0000_0422;
            12'o0103: crom <= 108'o3474_4751_1203_4374_4367_0700_0000_0000_0421;
            12'o0104: crom <= 108'o3676_3333_0004_7174_4007_0700_0410_0000_0212;
            12'o0105: crom <= 108'o0104_4751_1217_4374_4007_0700_0000_0000_0002;
            12'o0106: crom <= 108'o0110_4221_0011_4364_4277_0700_0200_0000_0010;
            12'o0107: crom <= 108'o0117_3443_0100_4174_4007_0700_0200_0014_0012;
            12'o0110: crom <= 108'o0125_4221_0010_4174_4477_0700_0000_0000_0000;
            12'o0111: crom <= 108'o3474_4751_1203_4374_4367_0700_0000_0000_0423;
            12'o0112: crom <= 108'o3474_4751_1203_4374_4367_0700_0000_0000_0422;
            12'o0113: crom <= 108'o3474_4751_1203_4374_4367_0700_0000_0000_0421;
            12'o0114: crom <= 108'o3675_4223_0000_4364_4277_0700_0210_0000_0010;
            12'o0115: crom <= 108'o0104_4751_1217_4374_4007_0700_0000_0000_0002;
            12'o0116: crom <= 108'o3674_4221_0004_4174_4007_0700_0200_0021_1016;
            12'o0117: crom <= 108'o0363_3771_0002_4365_5617_0700_0200_0000_0002;
            12'o0120: crom <= 108'o2774_4557_0006_1274_4007_0701_0010_0000_1441;
            12'o0121: crom <= 108'o2764_4557_0004_1274_4007_0701_0000_0000_1442;
            12'o0122: crom <= 108'o0122_3336_0604_4174_4046_2630_2000_0060_0000;
            12'o0123: crom <= 108'o0004_3334_0604_4174_4004_1700_0000_0000_0000;
            12'o0124: crom <= 108'o0171_3223_0000_1174_4007_0700_0400_0000_1443;
            12'o0125: crom <= 108'o0131_4221_0013_4174_4257_0700_0000_0000_0000;
            12'o0126: crom <= 108'o0142_1116_0604_4174_4046_2630_6000_0060_0000;
            12'o0127: crom <= 108'o0004_1114_0604_4174_4004_1700_4000_0000_0000;
            12'o0130: crom <= 108'o3075_3771_0003_0276_6007_0700_0010_0000_0000;
            12'o0131: crom <= 108'o0162_3333_0013_7174_4007_0700_0400_0000_0230;
            12'o0132: crom <= 108'o2055_4221_0017_4174_4007_0700_0010_0000_0000;
            12'o0133: crom <= 108'o2030_3441_0305_1174_4007_0421_0000_0000_1441;
            12'o0134: crom <= 108'o3671_3441_0104_4170_4007_0700_0010_0000_0000;
            12'o0135: crom <= 108'o1400_0551_0501_4370_4007_0701_0000_0000_0001;
            12'o0136: crom <= 108'o1400_4113_0305_4174_4007_0330_0000_0000_0020;
            12'o0137: crom <= 108'o3613_3771_0005_4374_0007_0700_0000_0003_0130;
            12'o0140: crom <= 108'o0104_4751_1217_4374_4007_0700_0000_0000_1005;
            12'o0141: crom <= 108'o3607_4221_0014_4174_4007_0700_0010_0000_0000;
            12'o0142: crom <= 108'o0122_0116_0604_4174_4046_2630_2000_0060_0000;
            12'o0143: crom <= 108'o0004_0114_0604_4174_4004_1700_0000_0000_0000;
            12'o0144: crom <= 108'o3043_4222_0000_4174_4007_0700_2010_0071_0033;
            12'o0145: crom <= 108'o0144_3447_0303_4174_4007_0700_1000_0041_0001;
            12'o0146: crom <= 108'o0142_3336_0604_4174_4046_2630_2000_0060_0000;
            12'o0147: crom <= 108'o0004_3334_0604_4174_4004_1700_0000_0000_0000;
            12'o0150: crom <= 108'o2551_3771_0002_4365_5217_0700_0210_0000_0002;
            12'o0151: crom <= 108'o0343_4751_1217_4374_4007_0700_0000_0000_0120;
            12'o0152: crom <= 108'o0110_3441_0301_4170_4156_4700_0200_0014_0012;
            12'o0153: crom <= 108'o2055_3444_1616_4174_4067_0700_0010_0000_0000;
            12'o0154: crom <= 108'o3204_3227_0003_4174_4007_0700_0000_0000_0000;
            12'o0155: crom <= 108'o2054_3333_0003_4174_4007_0621_0010_0000_0000;
            12'o0156: crom <= 108'o2054_3333_0003_4174_4007_0621_0010_0000_0000;
            12'o0157: crom <= 108'o3204_3227_0003_4174_4007_0700_0000_0000_0000;
            12'o0160: crom <= 108'o1216_7443_0300_4174_4007_0621_0000_0000_0000;
            12'o0161: crom <= 108'o0164_3333_0005_4174_4007_0621_0000_0000_0000;
            12'o0162: crom <= 108'o0212_3333_0013_7174_4007_0700_0400_0000_0300;
            12'o0163: crom <= 108'o3000_3446_0606_4174_4007_0700_0010_0000_0000;
            12'o0164: crom <= 108'o0370_4443_0000_4174_4007_0700_2010_0071_0042;
            12'o0165: crom <= 108'o0555_4443_0000_4174_4467_0700_0000_0051_1000;
            12'o0166: crom <= 108'o1177_3441_0304_4174_4007_0700_0000_0000_0000;
            12'o0167: crom <= 108'o3177_4662_0000_4370_4007_0700_0000_0077_7000;
            12'o0170: crom <= 108'o0172_0551_0505_2270_4007_0700_0000_0000_0000;
            12'o0171: crom <= 108'o0563_3442_0300_4174_4007_0700_2010_0071_0043;
            12'o0172: crom <= 108'o0556_5741_0505_4174_4003_7700_0200_0000_0010;
            12'o0173: crom <= 108'o3225_3444_1616_4174_4067_0700_0000_0000_0000;
            12'o0174: crom <= 108'o3263_0551_0505_2270_4007_0700_0200_0004_0512;
            12'o0175: crom <= 108'o2763_3441_0416_4174_4007_0700_0000_0000_0000;
            12'o0176: crom <= 108'o3263_3443_0500_4174_4007_0700_0200_0004_0512;
            12'o0177: crom <= 108'o3204_2227_0003_4174_4007_0700_4000_0000_0000;
            12'o0200: crom <= 108'o0200_3444_0303_4174_4043_4701_1000_0041_1777;
            12'o0201: crom <= 108'o0110_0551_0201_2270_4156_4700_0200_0014_0012;
            12'o0202: crom <= 108'o0322_3333_0003_4174_4003_4701_0010_0000_0000;
            12'o0203: crom <= 108'o0110_3441_0201_4170_4156_4700_0200_0014_0012;
            12'o0204: crom <= 108'o0322_3446_0303_4174_4047_0700_1010_0041_0001;
            12'o0205: crom <= 108'o0366_0551_0202_2270_4007_0700_0200_0004_0012;
            12'o0206: crom <= 108'o0322_3446_0303_4174_4047_0700_1010_0041_0001;
            12'o0207: crom <= 108'o0366_3443_0200_4174_4007_0700_0200_0004_0012;
            12'o0210: crom <= 108'o3255_4002_0000_4174_0007_0700_0000_0000_0000;
            12'o0211: crom <= 108'o0213_0551_0202_2270_4007_0700_0000_0000_0000;
            12'o0212: crom <= 108'o0214_3333_0013_7174_4007_0700_0400_0000_0301;
            12'o0213: crom <= 108'o0000_5741_0203_4174_4001_3700_0200_0000_0342;
            12'o0214: crom <= 108'o0223_4223_0000_1174_4007_0700_0400_0000_1443;
            12'o0215: crom <= 108'o0366_0551_0202_2270_4007_0700_0200_0004_0112;
            12'o0216: crom <= 108'o0610_4111_1204_4174_4007_0700_0000_0000_0000;
            12'o0217: crom <= 108'o0366_3443_0200_4174_4007_0700_0200_0004_0112;
            12'o0220: crom <= 108'o0221_3441_0301_4174_4007_0700_0200_0014_0012;
            12'o0221: crom <= 108'o0100_3440_0404_0174_4156_4700_0400_0000_0000;
            12'o0222: crom <= 108'o1400_3440_0404_0174_4007_0700_0400_0000_0000;
            12'o0223: crom <= 108'o0226_3333_0007_1174_4007_0700_0400_0000_1444;
            12'o0224: crom <= 108'o0323_4443_0000_4174_4007_0700_0000_0000_0000;
            12'o0225: crom <= 108'o0140_6553_0500_4374_4007_0321_0000_0033_0656;
            12'o0226: crom <= 108'o0235_4221_0003_4174_4007_0700_2000_0071_0023;
            12'o0227: crom <= 108'o2452_4553_0300_4374_4007_0331_0000_0000_0001;
            12'o0230: crom <= 108'o3101_0553_0300_2274_4007_0701_0200_0004_0712;
            12'o0231: crom <= 108'o3447_3441_0503_4174_4007_0700_0000_0000_0000;
            12'o0232: crom <= 108'o3101_3443_0300_4174_4007_0700_0200_0004_0712;
            12'o0233: crom <= 108'o3446_3770_0503_4334_4017_0700_0000_0032_6000;
            12'o0234: crom <= 108'o3454_0553_0300_2274_4007_0701_0200_0004_0612;
            12'o0235: crom <= 108'o0242_3333_0007_7174_4007_0700_0400_0000_0344;
            12'o0236: crom <= 108'o3454_3443_0300_4174_4007_0700_0200_0004_0612;
            12'o0237: crom <= 108'o3650_4571_1204_4374_4007_0700_0000_0021_1200;
            12'o0240: crom <= 108'o3127_3333_0003_7174_4007_0700_0400_0000_0223;
            12'o0241: crom <= 108'o0350_3770_0305_4334_4016_7351_0010_0033_6000;
            12'o0242: crom <= 108'o0244_4223_0000_7174_4007_0700_0400_0000_0373;
            12'o0243: crom <= 108'o2054_3333_0017_4174_4007_0621_0010_0000_0000;
            12'o0244: crom <= 108'o0311_3771_0002_4374_4007_0700_0000_0000_0344;
            12'o0245: crom <= 108'o0110_3443_0100_4174_4156_4700_0200_0014_0012;
            12'o0246: crom <= 108'o3412_3333_0004_7174_4007_0700_0410_0000_0246;
            12'o0247: crom <= 108'o3411_3771_0003_7274_4007_0701_0000_0000_0246;
            12'o0250: crom <= 108'o0110_3443_0100_4174_4156_4700_0200_0014_0012;
            12'o0251: crom <= 108'o1400_3333_0003_4174_4007_0520_0000_0000_0000;
            12'o0252: crom <= 108'o1400_3333_0003_4174_4007_0621_0000_0000_0000;
            12'o0253: crom <= 108'o1400_3333_0003_4174_4007_0421_0000_0000_0000;
            12'o0254: crom <= 108'o0110_0111_0701_4170_4156_4700_0200_0014_0012;
            12'o0255: crom <= 108'o0260_3333_0003_4174_4007_0520_0000_0000_0000;
            12'o0256: crom <= 108'o0260_3333_0003_4174_4007_0621_0000_0000_0000;
            12'o0257: crom <= 108'o0260_3333_0003_4174_4007_0421_0000_0000_0000;
            12'o0260: crom <= 108'o0110_0111_0701_4170_4156_4700_0200_0014_0012;
            12'o0261: crom <= 108'o0110_3443_0100_4174_4156_4700_0200_0014_0012;
            12'o0262: crom <= 108'o0407_3447_0705_4174_4003_7700_0000_0000_0000;
            12'o0263: crom <= 108'o3236_3444_0303_4174_4047_0700_0000_0000_0000;
            12'o0264: crom <= 108'o3077_3333_0003_4174_4217_0700_0010_0000_0500;
            12'o0265: crom <= 108'o0360_3333_0003_4174_4006_5701_0010_0000_0000;
            12'o0266: crom <= 108'o0262_3447_0303_4174_4007_0700_1000_0041_0001;
            12'o0267: crom <= 108'o1400_4443_0000_4174_4467_0700_0000_0005_0000;
            12'o0270: crom <= 108'o0100_3440_0505_0174_4156_4700_0400_0000_0000;
            12'o0271: crom <= 108'o0762_3770_0505_0174_4007_0520_0400_0000_0000;
            12'o0272: crom <= 108'o0762_3770_0505_0174_4007_0621_0400_0000_0000;
            12'o0273: crom <= 108'o0762_3770_0505_0174_4007_0421_0400_0000_0000;
            12'o0274: crom <= 108'o0764_3440_0505_0174_4007_0700_0400_0000_0000;
            12'o0275: crom <= 108'o0764_3770_0505_0174_4007_0520_0400_0000_0000;
            12'o0276: crom <= 108'o0764_3770_0505_0174_4007_0621_0400_0000_0000;
            12'o0277: crom <= 108'o0764_3770_0505_0174_4007_0421_0400_0000_0000;
            12'o0300: crom <= 108'o2737_4551_0202_4374_0007_0700_0000_0077_7740;
            12'o0301: crom <= 108'o2551_3771_0002_4365_5217_0700_0210_0000_0002;
            12'o0302: crom <= 108'o0016_4443_0000_4174_4004_1700_0000_0000_0000;
            12'o0303: crom <= 108'o2432_4553_1400_4374_4007_0331_0010_0007_7400;
            12'o0304: crom <= 108'o0305_5111_0514_4170_4007_0700_0000_0000_0000;
            12'o0305: crom <= 108'o3610_3770_1416_4344_4007_0700_0010_0000_0000;
            12'o0306: crom <= 108'o0016_3447_0303_4174_4004_1700_1000_0041_0001;
            12'o0307: crom <= 108'o3610_3770_1416_4344_4007_0700_0010_0000_0000;
            12'o0310: crom <= 108'o2746_3333_0002_4175_5007_0701_0210_0000_0002;
            12'o0311: crom <= 108'o0323_3771_0006_4374_4007_0700_0000_0000_0373;
            12'o0312: crom <= 108'o2745_3741_0103_4074_4007_0700_0010_0000_0000;
            12'o0313: crom <= 108'o0022_3333_0003_4175_5007_0701_0200_0000_0002;
            12'o0314: crom <= 108'o2746_3333_0003_4175_5007_0701_0210_0000_0002;
            12'o0315: crom <= 108'o0110_3443_0100_4174_4156_4700_0200_0014_0012;
            12'o0316: crom <= 108'o0020_3333_0001_4175_5007_0701_0200_0000_0002;
            12'o0317: crom <= 108'o0110_3441_0301_4170_4156_4700_0200_0014_0012;
            12'o0320: crom <= 108'o2737_4551_0202_4374_0007_0700_0000_0077_7740;
            12'o0321: crom <= 108'o2432_4553_1400_4374_4007_0331_0010_0007_7400;
            12'o0322: crom <= 108'o0462_0007_0704_4174_4007_0511_0000_0000_0000;
            12'o0323: crom <= 108'o0010_0111_0706_4174_4007_0700_0200_0000_0010;
            12'o0324: crom <= 108'o0334_0111_0702_4174_4007_0700_0200_0000_0010;
            12'o0325: crom <= 108'o0335_3333_0012_4174_4437_0700_0000_0000_0000;
            12'o0326: crom <= 108'o0322_3446_0303_4174_4047_0700_1000_0041_0001;
            12'o0327: crom <= 108'o2002_4553_1300_4374_4007_0321_0000_0000_2000;
            12'o0330: crom <= 108'o1220_3333_0005_4174_4007_0520_0000_0000_0000;
            12'o0331: crom <= 108'o3071_4551_0404_4374_0007_0700_0010_0037_7777;
            12'o0332: crom <= 108'o3450_3771_0003_7274_4007_0700_0010_0000_0244;
            12'o0333: crom <= 108'o1220_3333_0005_4174_4007_0520_0000_0000_0000;
            12'o0334: crom <= 108'o0224_3333_0004_6174_4007_0630_2400_0060_0000;
            12'o0335: crom <= 108'o1525_4223_0000_4364_4277_0700_0200_0000_0010;
            12'o0336: crom <= 108'o3437_3771_0003_1276_6007_0701_0000_0000_1443;
            12'o0337: crom <= 108'o2005_4111_1203_4174_4007_0700_0000_0000_0000;
            12'o0340: crom <= 108'o0550_4443_0000_4174_4006_7701_0000_0031_0210;
            12'o0341: crom <= 108'o3102_3770_0505_4334_4057_0700_0000_0073_0000;
            12'o0342: crom <= 108'o3102_3770_0505_4334_4057_0700_0000_0074_0000;
            12'o0343: crom <= 108'o0346_4221_0001_4174_4467_0700_0000_0000_0004;
            12'o0344: crom <= 108'o3102_3770_0505_4334_4057_0700_0000_0075_0000;
            12'o0345: crom <= 108'o3102_3770_0505_4334_4057_0700_0000_0076_0000;
            12'o0346: crom <= 108'o0116_3771_0017_4374_4007_0700_0000_0000_0000;
            12'o0347: crom <= 108'o3102_3770_0505_4334_4057_0700_0000_0077_0000;
            12'o0350: crom <= 108'o3075_3441_0503_4174_4007_0700_0200_0003_0002;
            12'o0351: crom <= 108'o0004_4443_0000_4174_4004_1700_0000_0000_0000;
            12'o0352: crom <= 108'o3074_3770_0503_4334_4017_0700_0000_0032_6000;
            12'o0353: crom <= 108'o0004_4443_0000_4174_4004_1700_0000_0000_0000;
            12'o0354: crom <= 108'o1264_3446_1200_4174_4007_0700_2010_0071_0042;
            12'o0355: crom <= 108'o3040_3444_0303_4174_4047_0700_0000_0000_0000;
            12'o0356: crom <= 108'o3021_3224_0016_4174_4007_0700_0000_0000_0000;
            12'o0357: crom <= 108'o3037_2222_0000_4174_4007_0700_4000_0000_0000;
            12'o0360: crom <= 108'o3114_3333_0003_4174_4007_0700_1000_0031_7770;
            12'o0361: crom <= 108'o3112_3770_0503_4334_4017_0700_0000_0041_0000;
            12'o0362: crom <= 108'o3112_3770_0503_4334_4027_0700_0000_0041_0000;
            12'o0363: crom <= 108'o0201_0111_0701_2170_4366_6700_0200_0010_0010;
            12'o0364: crom <= 108'o3112_3770_0503_4334_4037_0700_0000_0041_0000;
            12'o0365: crom <= 108'o3112_3770_0503_4334_4047_0700_0000_0041_0000;
            12'o0366: crom <= 108'o0371_3771_0002_4361_5217_0700_0200_0000_0102;
            12'o0367: crom <= 108'o3112_3770_0503_4334_4057_0700_0000_0041_0000;
            12'o0370: crom <= 108'o3043_4662_0000_4374_0007_0700_0010_0037_7777;
            12'o0371: crom <= 108'o0201_3443_0100_2174_4006_6700_0200_0010_0010;
            12'o0372: crom <= 108'o0412_3333_0003_4174_4007_0520_3010_0041_2000;
            12'o0373: crom <= 108'o0000_4221_0004_4174_4001_2700_0000_0000_0000;
            12'o0374: crom <= 108'o0002_4443_0000_4174_4004_1700_0000_0000_0000;
            12'o0375: crom <= 108'o0002_2222_0000_4174_4004_1700_4000_0000_0000;
            12'o0376: crom <= 108'o0377_2222_0000_4174_4007_0700_4000_0000_0000;
            12'o0377: crom <= 108'o0002_2441_0303_4174_4004_1700_4000_0000_0000;
            12'o0400: crom <= 108'o2747_3333_0003_4174_4007_0700_0200_0003_0012;
            12'o0401: crom <= 108'o0406_0111_0702_4170_4007_0700_0200_0004_0312;
            12'o0402: crom <= 108'o0445_0111_0703_4174_4007_0700_0200_0004_0312;
            12'o0403: crom <= 108'o0432_0111_0703_4174_4007_0700_0200_0004_0312;
            12'o0404: crom <= 108'o2737_4551_0202_4374_0007_0700_0000_0077_7740;
            12'o0405: crom <= 108'o0000_4443_0000_4174_4001_2700_0000_0000_0000;
            12'o0406: crom <= 108'o0000_3771_0004_4365_5001_2700_0200_0000_0002;
            12'o0407: crom <= 108'o0016_4443_0000_4174_4004_1700_0000_0000_0000;
            12'o0410: crom <= 108'o2775_3777_0006_0274_4007_0701_0010_0000_0000;
            12'o0411: crom <= 108'o2777_0113_1616_1174_4007_0701_0400_0000_1441;
            12'o0412: crom <= 108'o0001_4551_0303_4374_0004_1700_0000_0000_0777;
            12'o0413: crom <= 108'o0001_3551_0303_4374_0004_1700_0000_0077_7000;
            12'o0414: crom <= 108'o2765_3223_0000_1174_4007_0700_0400_0000_1442;
            12'o0415: crom <= 108'o0000_3771_0004_1276_6001_2701_0000_0000_1441;
            12'o0416: crom <= 108'o0431_3776_0005_0274_4007_0701_0000_0000_0000;
            12'o0417: crom <= 108'o0302_0111_0503_4174_4003_4701_0000_0000_0000;
            12'o0420: crom <= 108'o0420_3444_0303_4174_4063_4701_1000_0041_1777;
            12'o0421: crom <= 108'o2000_2222_0000_4174_4007_0311_4000_0000_0000;
            12'o0422: crom <= 108'o0262_3333_0003_4174_4003_4701_0010_0000_0000;
            12'o0423: crom <= 108'o2000_2222_0000_4174_4007_0311_4000_0000_0000;
            12'o0424: crom <= 108'o0262_3447_0303_4174_4007_0700_1010_0041_0001;
            12'o0425: crom <= 108'o2000_2222_0000_4174_4007_0311_4000_0000_0000;
            12'o0426: crom <= 108'o0262_3447_0303_4174_4007_0700_1010_0041_0001;
            12'o0427: crom <= 108'o2000_2222_0000_4174_4007_0311_4000_0000_0000;
            12'o0430: crom <= 108'o1376_3223_0000_4174_4007_0621_0000_0000_0000;
            12'o0431: crom <= 108'o0044_3446_0505_4174_4007_0700_0000_0000_0000;
            12'o0432: crom <= 108'o0451_3551_0505_4374_0007_0700_0000_0077_7000;
            12'o0433: crom <= 108'o3222_5111_1217_4174_4007_0700_0000_0000_0000;
            12'o0434: crom <= 108'o1515_3333_0003_4175_5007_0701_0200_0000_0002;
            12'o0435: crom <= 108'o1400_3333_0003_4175_5007_0701_0200_0000_0002;
            12'o0436: crom <= 108'o1377_3770_0303_4324_0457_0700_0000_0041_0000;
            12'o0437: crom <= 108'o0433_0222_0000_4174_4007_0700_4000_0000_0000;
            12'o0440: crom <= 108'o0440_3444_0303_4174_4063_4701_1000_0041_1777;
            12'o0441: crom <= 108'o2214_3771_0004_1276_6007_0701_0010_0000_1441;
            12'o0442: crom <= 108'o0262_3333_0003_4174_4003_4701_0010_0000_0000;
            12'o0443: crom <= 108'o2170_0111_0706_4174_4007_0630_2000_0060_0000;
            12'o0444: crom <= 108'o0262_3447_0303_4174_4007_0700_1010_0041_0001;
            12'o0445: crom <= 108'o0451_4551_0505_4374_0007_0700_0000_0000_0777;
            12'o0446: crom <= 108'o0262_3447_0303_4174_4007_0700_1010_0041_0001;
            12'o0447: crom <= 108'o2172_4553_0600_4374_4007_0331_0000_0077_7777;
            12'o0450: crom <= 108'o0440_3444_0303_4174_4063_4701_1000_0041_1777;
            12'o0451: crom <= 108'o0452_4557_0004_4365_5007_0701_0200_0000_0002;
            12'o0452: crom <= 108'o0467_3447_0503_4174_4007_0700_0000_0000_0000;
            12'o0453: crom <= 108'o3227_3446_1616_4174_4047_0700_0000_0000_0000;
            12'o0454: crom <= 108'o0454_3444_0303_4174_4447_0630_2000_0060_0000;
            12'o0455: crom <= 108'o1515_3445_0303_4174_4007_0700_0000_0000_0000;
            12'o0456: crom <= 108'o0327_3770_0303_4324_0453_7700_0000_0041_0000;
            12'o0457: crom <= 108'o0453_3551_1313_4374_0007_0700_0000_0000_2000;
            12'o0460: crom <= 108'o1074_0551_0703_7274_4007_0701_0010_0000_0242;
            12'o0461: crom <= 108'o2142_4553_0600_4374_4007_0321_0000_0010_0000;
            12'o0462: crom <= 108'o0016_3770_0303_4324_0454_1700_0000_0041_0000;
            12'o0463: crom <= 108'o0462_0441_0303_4174_4003_4701_4000_0000_0000;
            12'o0464: crom <= 108'o3335_7771_0003_7274_4007_0701_0000_0000_0242;
            12'o0465: crom <= 108'o2132_1553_0300_4374_4007_0532_4000_0000_0012;
            12'o0466: crom <= 108'o0462_3447_0303_4174_4007_0700_1000_0041_0001;
            12'o0467: crom <= 108'o0471_3447_0303_4174_4007_0700_2000_0011_0000;
            12'o0470: crom <= 108'o3667_3741_0105_4074_4007_0700_0010_0000_0000;
            12'o0471: crom <= 108'o0000_3443_0100_4174_4001_2700_0200_0014_0012;
            12'o0472: crom <= 108'o0472_3446_1616_4174_4046_2630_2000_0060_0000;
            12'o0473: crom <= 108'o0453_3221_0017_4174_4006_2700_0000_0000_0000;
            12'o0474: crom <= 108'o3664_3771_0003_4374_0007_0700_0010_0000_0000;
            12'o0475: crom <= 108'o2714_3441_0301_4174_4467_0700_0000_0000_0004;
            12'o0476: crom <= 108'o2016_3551_1313_4374_0007_0700_0000_0000_2000;
            12'o0477: crom <= 108'o2017_3551_1313_4374_0007_0700_0000_0000_2000;
            12'o0500: crom <= 108'o1074_0551_0703_7274_4007_0701_0010_0000_0242;
            12'o0501: crom <= 108'o0750_3441_0304_4174_4007_0520_0000_0000_0000;
            12'o0502: crom <= 108'o0767_3441_0301_4174_4007_0700_0200_0014_0012;
            12'o0503: crom <= 108'o1400_4223_0000_1174_4007_0700_0400_0000_1441;
            12'o0504: crom <= 108'o3270_1771_0003_7274_4007_0701_4000_0000_0242;
            12'o0505: crom <= 108'o3450_3771_0013_4370_4007_0700_0010_0000_0005;
            12'o0506: crom <= 108'o1515_3333_0005_4175_5007_0701_0200_0000_0002;
            12'o0507: crom <= 108'o0500_3771_0013_4370_4007_0700_0000_0000_0003;
            12'o0510: crom <= 108'o3450_3771_0013_4370_4007_0700_0010_0000_0012;
            12'o0511: crom <= 108'o1402_3771_0003_0270_6007_0700_0000_0000_0000;
            12'o0512: crom <= 108'o1402_3771_0003_0276_0007_0700_0000_0000_0000;
            12'o0513: crom <= 108'o2040_3333_0017_4174_4007_0520_1000_0031_0202;
            12'o0514: crom <= 108'o0514_3445_0505_4174_4007_0520_1000_0041_0004;
            12'o0515: crom <= 108'o1006_3777_0003_4334_4057_0700_0000_0041_0000;
            12'o0516: crom <= 108'o3365_2551_0705_1274_4007_0701_4000_0000_1443;
            12'o0517: crom <= 108'o0513_0222_0000_4174_4007_0700_4000_0000_0000;
            12'o0520: crom <= 108'o0520_3444_0303_4174_4043_4701_1000_0041_1777;
            12'o0521: crom <= 108'o2044_4553_1300_4374_4007_0321_0000_0000_2000;
            12'o0522: crom <= 108'o0322_3333_0003_4174_4003_4701_0010_0000_0000;
            12'o0523: crom <= 108'o2044_4553_1300_4374_4007_0321_0000_0000_2000;
            12'o0524: crom <= 108'o0322_3446_0303_4174_4047_0700_1010_0041_0001;
            12'o0525: crom <= 108'o2044_4553_1300_4374_4007_0321_0000_0000_2000;
            12'o0526: crom <= 108'o0322_3446_0303_4174_4047_0700_1010_0041_0001;
            12'o0527: crom <= 108'o2044_4553_1300_4374_4007_0321_0000_0000_2000;
            12'o0530: crom <= 108'o3251_4002_0000_4174_0007_0700_0000_0000_0000;
            12'o0531: crom <= 108'o0532_3333_0004_4175_5007_0701_0200_0000_0002;
            12'o0532: crom <= 108'o0435_3443_0200_4174_4007_0700_0200_0003_0312;
            12'o0533: crom <= 108'o3444_1111_0703_4174_4007_0700_4000_0000_0000;
            12'o0534: crom <= 108'o0534_3446_0505_4174_4057_0630_2000_0060_0000;
            12'o0535: crom <= 108'o1033_3444_0505_4174_4007_0700_0000_0000_0000;
            12'o0536: crom <= 108'o3250_4221_0013_4174_4007_0700_0000_0000_0000;
            12'o0537: crom <= 108'o1074_0551_0703_7274_4007_0701_0000_0000_0242;
            12'o0540: crom <= 108'o2274_3333_0004_7174_4007_0520_0410_0000_0242;
            12'o0541: crom <= 108'o0750_3441_0304_4174_4007_0520_0000_0000_0000;
            12'o0542: crom <= 108'o3450_3771_0013_4370_4007_0700_0010_0000_0005;
            12'o0543: crom <= 108'o0563_3442_0300_4174_4007_0700_2010_0071_0043;
            12'o0544: crom <= 108'o0544_3444_0505_4174_4057_0630_2000_0060_0000;
            12'o0545: crom <= 108'o1033_3444_0505_4174_4007_0700_0000_0000_0000;
            12'o0546: crom <= 108'o3306_0551_0704_7274_4007_0701_0000_0000_0242;
            12'o0547: crom <= 108'o2766_3445_0404_4174_4467_0700_0000_0005_0000;
            12'o0550: crom <= 108'o3104_4443_0000_4174_4007_0700_1000_0031_0000;
            12'o0551: crom <= 108'o1264_3446_0316_4174_4007_0520_2010_0071_0042;
            12'o0552: crom <= 108'o3103_3770_0505_4344_4007_0700_0000_0000_0000;
            12'o0553: crom <= 108'o3024_3224_0016_4174_4007_0700_0000_0000_0000;
            12'o0554: crom <= 108'o1046_3772_0000_1275_5007_0701_0000_0000_1441;
            12'o0555: crom <= 108'o0100_4443_0000_4174_4156_4700_0000_0000_0000;
            12'o0556: crom <= 108'o3400_3333_0005_7174_4001_2700_0400_0000_0241;
            12'o0557: crom <= 108'o2056_3333_0005_4174_4007_0530_0000_0000_0000;
            12'o0560: crom <= 108'o0620_3771_0005_1276_6007_0701_0010_0000_1443;
            12'o0561: crom <= 108'o2140_0551_0404_1274_4007_0562_0010_0000_1444;
            12'o0562: crom <= 108'o2214_0111_0705_4174_4007_0700_0010_0000_0000;
            12'o0563: crom <= 108'o3002_3446_1200_4174_4007_0700_0010_0000_0000;
            12'o0564: crom <= 108'o1500_3111_0503_4174_4003_7700_0200_0003_0001;
            12'o0565: crom <= 108'o0600_0551_0505_1274_4007_0701_0000_0000_1443;
            12'o0566: crom <= 108'o3364_3333_0003_7174_4007_0700_0400_0000_0247;
            12'o0567: crom <= 108'o0004_0113_0404_4174_4464_1701_0000_0001_0001;
            12'o0570: crom <= 108'o0571_3771_0003_4374_4007_0700_0000_0000_0000;
            12'o0571: crom <= 108'o0370_3333_0005_7174_4007_0700_0410_0000_0226;
            12'o0572: crom <= 108'o1515_3445_0303_4174_4007_0700_1020_0041_0001;
            12'o0573: crom <= 108'o3143_3772_0000_4374_0007_0700_0000_0000_0000;
            12'o0574: crom <= 108'o0500_3771_0013_4370_4007_0700_0000_0000_0003;
            12'o0575: crom <= 108'o3265_3771_0005_1276_6007_0701_0000_0000_1444;
            12'o0576: crom <= 108'o3305_3441_0304_4174_4007_0700_0000_0000_0000;
            12'o0577: crom <= 108'o0630_3771_0004_1276_6007_0522_0000_0000_1443;
            12'o0600: crom <= 108'o0621_4443_0000_4174_4007_0700_0010_0000_0000;
            12'o0601: crom <= 108'o2140_0111_0304_4174_4007_0561_0010_0000_0000;
            12'o0602: crom <= 108'o0602_3445_0303_4174_4007_0630_2000_0060_0000;
            12'o0603: crom <= 108'o3772_4443_0000_4174_4007_0700_0010_0000_0000;
            12'o0604: crom <= 108'o0340_3333_0003_4174_4006_5701_1010_0051_0770;
            12'o0605: crom <= 108'o3333_3440_0404_1174_4007_0700_0400_0000_1444;
            12'o0606: crom <= 108'o0555_3440_0303_0174_4467_0700_0400_0005_0000;
            12'o0607: crom <= 108'o1000_4443_0000_4174_4007_0700_0000_0000_0000;
            12'o0610: crom <= 108'o3256_4111_0004_4174_4007_0700_0010_0000_0000;
            12'o0611: crom <= 108'o1515_3447_0303_4174_4007_0700_1020_0041_0001;
            12'o0612: crom <= 108'o3253_6111_0004_4174_4007_0700_0000_0000_0000;
            12'o0613: crom <= 108'o2050_2441_0404_4174_4007_0561_4000_0000_0000;
            12'o0614: crom <= 108'o0634_3447_0505_4174_4007_0700_2000_0041_1776;
            12'o0615: crom <= 108'o0624_3447_0505_4174_4007_0700_2000_0031_1776;
            12'o0616: crom <= 108'o3330_3771_0013_4370_4007_0700_0000_0000_0007;
            12'o0617: crom <= 108'o0616_3551_0606_4374_0007_0700_0000_0040_0000;
            12'o0620: crom <= 108'o0621_4443_0000_4174_4007_0700_0010_0000_0000;
            12'o0621: crom <= 108'o0622_0111_0505_4174_4007_0700_0000_0000_0000;
            12'o0622: crom <= 108'o2140_0111_0404_4174_4007_0561_0010_0000_0000;
            12'o0623: crom <= 108'o3001_3447_0606_4174_4007_0700_2010_0071_0043;
            12'o0624: crom <= 108'o0624_3446_0505_4174_4047_0630_2000_0060_0000;
            12'o0625: crom <= 108'o1053_3444_0505_4174_4047_0700_0000_0000_0000;
            12'o0626: crom <= 108'o0001_4443_0000_4174_4004_1700_0000_0000_0000;
            12'o0627: crom <= 108'o0730_3442_0300_4174_4007_0700_2000_0071_0043;
            12'o0630: crom <= 108'o3274_3771_0003_1276_6007_0701_0000_0000_1441;
            12'o0631: crom <= 108'o2263_3771_0013_4370_4007_0700_0010_0000_0006;
            12'o0632: crom <= 108'o0454_3777_0003_0274_4007_0631_2000_0060_0000;
            12'o0633: crom <= 108'o3306_0551_0704_7274_4007_0701_0000_0000_0242;
            12'o0634: crom <= 108'o0634_3444_0505_4174_4447_0630_2000_0060_0000;
            12'o0635: crom <= 108'o1053_3444_0505_4174_4447_0700_0000_0000_0000;
            12'o0636: crom <= 108'o2206_3333_0003_4174_4007_0700_0200_0004_0012;
            12'o0637: crom <= 108'o0510_3333_0004_7174_4007_0700_0400_0000_0250;
            12'o0640: crom <= 108'o2157_3440_0606_1174_4007_0700_0400_0000_1443;
            12'o0641: crom <= 108'o3450_3333_0005_7174_4007_0700_0410_0000_0242;
            12'o0642: crom <= 108'o1064_4662_0000_4374_0007_0700_0000_0037_7777;
            12'o0643: crom <= 108'o1064_3662_0000_4374_0007_0700_0000_0040_0000;
            12'o0644: crom <= 108'o0644_3446_0505_4174_4077_0630_2000_0060_0000;
            12'o0645: crom <= 108'o1033_3444_0505_4174_4007_0700_0000_0000_0000;
            12'o0646: crom <= 108'o0701_3447_0303_4174_4007_0700_0000_0000_0000;
            12'o0647: crom <= 108'o3362_2551_0705_1274_4007_0701_4000_0000_1443;
            12'o0650: crom <= 108'o3274_3441_0503_4174_4007_0700_0000_0000_0000;
            12'o0651: crom <= 108'o3275_7771_0003_7274_4007_0701_0000_0000_0242;
            12'o0652: crom <= 108'o3276_3770_0503_4334_4017_0700_0000_0032_6000;
            12'o0653: crom <= 108'o3275_7771_0003_7274_4007_0701_0000_0000_0242;
            12'o0654: crom <= 108'o2226_3770_0303_4344_4007_0700_2000_0071_0007;
            12'o0655: crom <= 108'o2227_3770_0303_4344_4007_0700_0000_0000_0000;
            12'o0656: crom <= 108'o2226_3447_0303_4174_4007_0700_2000_0071_0006;
            12'o0657: crom <= 108'o3403_4551_0303_4374_4007_0700_0000_0000_0777;
            12'o0660: crom <= 108'o0370_3771_0003_4374_4007_0700_0010_0000_0000;
            12'o0661: crom <= 108'o2232_1553_0300_4374_4007_0532_4000_0000_0005;
            12'o0662: crom <= 108'o3135_3223_0000_7174_4007_0700_0400_0000_0224;
            12'o0663: crom <= 108'o2250_3333_0006_4174_4007_0520_0000_0000_0000;
            12'o0664: crom <= 108'o0370_3771_0003_4374_4007_0700_0010_0000_0000;
            12'o0665: crom <= 108'o3423_4443_0000_4174_4007_0700_0000_0000_0000;
            12'o0666: crom <= 108'o3141_3333_0003_7174_4007_0700_0400_0000_0225;
            12'o0667: crom <= 108'o3423_4443_0000_4174_4007_0700_0000_0000_0000;
            12'o0670: crom <= 108'o1334_3333_0005_4174_4007_0520_0000_0000_0000;
            12'o0671: crom <= 108'o3423_4443_0000_4174_4007_0700_0000_0000_0000;
            12'o0672: crom <= 108'o3172_3441_0304_4174_4007_0700_0000_0000_0000;
            12'o0673: crom <= 108'o2254_4553_0600_4374_4007_0321_0000_0010_0000;
            12'o0674: crom <= 108'o0555_4443_0000_4174_4467_0700_0000_0041_1000;
            12'o0675: crom <= 108'o2254_4553_0600_4374_4007_0321_0000_0020_0000;
            12'o0676: crom <= 108'o0720_4443_0000_4174_4006_7701_2000_0041_1544;
            12'o0677: crom <= 108'o2254_4443_0000_4174_4007_0700_0000_0000_0000;
            12'o0700: crom <= 108'o3443_0551_0303_7274_4007_0700_0010_0000_0241;
            12'o0701: crom <= 108'o0706_3447_0303_4174_4037_0700_1020_0041_0001;
            12'o0702: crom <= 108'o2244_3333_0003_4174_4007_0621_0000_0000_0000;
            12'o0703: crom <= 108'o0246_3771_0013_4370_4007_0700_0000_0000_0011;
            12'o0704: crom <= 108'o3404_4443_0000_4174_4007_0700_0000_0000_0000;
            12'o0705: crom <= 108'o3450_3771_0013_4370_4007_0700_0010_0000_0013;
            12'o0706: crom <= 108'o0455_3445_0303_4174_4007_0700_0000_0000_0000;
            12'o0707: crom <= 108'o3423_4443_0000_4174_4007_0700_0000_0000_0000;
            12'o0710: crom <= 108'o3404_0111_0701_4174_4007_0700_0000_0000_0000;
            12'o0711: crom <= 108'o2240_3771_0013_4370_4007_0700_0000_0000_0011;
            12'o0712: crom <= 108'o0006_3333_0006_4174_4007_0520_0000_0000_0000;
            12'o0713: crom <= 108'o3423_4551_0606_4374_0007_0700_0000_0007_7777;
            12'o0714: crom <= 108'o0715_3771_0005_1276_6007_0701_0000_0000_1443;
            12'o0715: crom <= 108'o2236_3443_0500_4174_4007_0700_0200_0004_0012;
            12'o0716: crom <= 108'o3442_3447_0303_4174_4007_0700_0000_0000_0000;
            12'o0717: crom <= 108'o3440_3770_0303_7174_0007_0700_0000_0000_0241;
            12'o0720: crom <= 108'o1370_4443_0000_4174_4007_0630_2000_0060_0000;
            12'o0721: crom <= 108'o2270_3333_0006_4174_4007_0520_0000_0000_0000;
            12'o0722: crom <= 108'o3210_4443_0000_4174_4007_0700_2000_0031_0232;
            12'o0723: crom <= 108'o0004_4443_0000_4174_4004_1700_0000_0000_0000;
            12'o0724: crom <= 108'o1264_4222_0000_4174_4007_0700_2010_0071_0032;
            12'o0725: crom <= 108'o0721_5551_0606_4374_0007_0700_0000_0010_0000;
            12'o0726: crom <= 108'o1054_3221_0016_4174_4007_0700_2000_0071_0043;
            12'o0727: crom <= 108'o0721_3551_0606_4374_0007_0700_0000_0010_0000;
            12'o0730: crom <= 108'o3002_4443_0000_4174_4007_0700_0010_0000_0000;
            12'o0731: crom <= 108'o0721_3551_0606_4374_0007_0700_0000_0020_0000;
            12'o0732: crom <= 108'o3002_3442_0500_4174_4007_0700_2010_0071_0043;
            12'o0733: crom <= 108'o0004_3551_0606_4374_0004_1700_0000_0020_0000;
            12'o0734: crom <= 108'o3233_3441_0416_4174_4007_0700_0000_0000_0000;
            12'o0735: crom <= 108'o0731_5551_0606_4374_0007_0700_0000_0010_0000;
            12'o0736: crom <= 108'o3235_3221_0017_4174_4007_0700_0000_0000_0000;
            12'o0737: crom <= 108'o0721_3551_0606_4374_0007_0700_0000_0030_0000;
            12'o0740: crom <= 108'o3450_3551_1313_4370_4007_0700_0010_0000_0012;
            12'o0741: crom <= 108'o3416_3551_0606_4374_0007_0700_0000_0040_0000;
            12'o0742: crom <= 108'o0742_3444_0505_4174_4077_0630_2000_0060_0000;
            12'o0743: crom <= 108'o1033_3444_0505_4174_4007_0700_0000_0000_0000;
            12'o0744: crom <= 108'o0250_3440_0303_0174_4003_7700_0400_0000_0000;
            12'o0745: crom <= 108'o0250_4443_0000_4174_4003_7700_0000_0000_0000;
            12'o0746: crom <= 108'o3416_3551_0606_4374_0007_0700_0000_0040_0000;
            12'o0747: crom <= 108'o0752_3447_0303_4174_4007_0700_0000_0000_0000;
            12'o0750: crom <= 108'o3307_4223_0000_1174_4007_0700_0400_0000_1443;
            12'o0751: crom <= 108'o2263_3771_0013_4370_4007_0700_0010_0000_0004;
            12'o0752: crom <= 108'o0706_3445_0303_4174_4037_0700_1020_0041_0001;
            12'o0753: crom <= 108'o2147_3440_0606_0174_4007_0700_0400_0000_0000;
            12'o0754: crom <= 108'o0533_3771_0003_1276_6003_7701_0000_0000_1443;
            12'o0755: crom <= 108'o2271_3551_0606_4374_0007_0700_0000_0040_0000;
            12'o0756: crom <= 108'o0002_3771_0003_7274_4004_1701_0000_0000_0244;
            12'o0757: crom <= 108'o0003_3771_0003_1276_6004_1701_0000_0000_1444;
            12'o0760: crom <= 108'o3450_3771_0013_4370_4007_0700_0010_0000_0012;
            12'o0761: crom <= 108'o3423_4443_0000_4174_4007_0700_0000_0000_0000;
            12'o0762: crom <= 108'o0110_3443_0100_4174_4156_4700_0200_0014_0012;
            12'o0763: crom <= 108'o0110_3441_0301_4170_4156_4700_0200_0014_0012;
            12'o0764: crom <= 108'o0110_3441_0301_4170_4156_4700_0200_0014_0012;
            12'o0765: crom <= 108'o0110_3443_0100_4174_4156_4700_0200_0014_0012;
            12'o0766: crom <= 108'o3423_4443_0000_4174_4007_0700_0000_0000_0000;
            12'o0767: crom <= 108'o0514_4443_0000_4174_4007_0700_1000_0071_1764;
            12'o0770: crom <= 108'o0770_3773_0000_4074_4003_1701_0000_0000_0000;
            12'o0771: crom <= 108'o3622_3551_1414_4370_4007_0700_0000_0004_0000;
            12'o0772: crom <= 108'o3623_3551_1414_4370_4007_0700_0000_0002_0000;
            12'o0773: crom <= 108'o3624_3551_1414_4370_4007_0700_0000_0001_0000;
            12'o0774: crom <= 108'o3625_3551_1414_4370_4007_0700_0000_0000_4000;
            12'o0775: crom <= 108'o3626_3551_1414_4370_4007_0700_0000_0000_2000;
            12'o0776: crom <= 108'o3627_3551_1414_4370_4007_0700_0000_0000_1000;
            12'o0777: crom <= 108'o3630_3551_1414_4370_4007_0700_0000_0000_0400;
            12'o1000: crom <= 108'o3767_4443_0000_4174_4007_0700_2010_0071_0007;
            12'o1001: crom <= 108'o2552_4553_0300_4374_4007_0321_0000_0000_0077;
            12'o1002: crom <= 108'o2550_0551_0303_7274_4007_0701_0000_0000_0215;
            12'o1003: crom <= 108'o3772_0551_0303_7274_4007_0701_0010_0000_0215;
            12'o1004: crom <= 108'o2737_4551_0202_4374_0007_0700_0000_0077_7740;
            12'o1005: crom <= 108'o2601_3441_0301_4174_4007_0700_0000_0000_0000;
            12'o1006: crom <= 108'o1023_4251_0303_4374_4007_0700_0000_0000_0077;
            12'o1007: crom <= 108'o2546_4553_0300_4374_4007_0321_0000_0000_0077;
            12'o1010: crom <= 108'o2737_4551_0202_4374_0007_0700_0000_0077_7740;
            12'o1011: crom <= 108'o0303_4443_0000_4174_4007_0700_0000_0000_0000;
            12'o1012: crom <= 108'o3002_3442_0300_4174_4007_0700_2010_0071_0043;
            12'o1013: crom <= 108'o3647_3551_0505_0274_4007_0700_0000_0000_0000;
            12'o1014: crom <= 108'o2737_4551_0202_4374_0007_0700_0000_0077_7740;
            12'o1015: crom <= 108'o0060_4521_1205_4074_4007_0700_0000_0000_0000;
            12'o1016: crom <= 108'o0243_3446_0403_4174_4007_0700_1000_0041_1576;
            12'o1017: crom <= 108'o3647_5551_0505_0274_4007_0700_0000_0000_0000;
            12'o1020: crom <= 108'o2275_3771_0013_4370_4007_0700_0010_0000_0011;
            12'o1021: crom <= 108'o2120_3333_0004_4174_4007_0520_0000_0000_0000;
            12'o1022: crom <= 108'o3312_3333_0003_7174_4007_0700_0400_0000_0245;
            12'o1023: crom <= 108'o0100_3440_0303_1174_4156_4700_0400_0000_1441;
            12'o1024: crom <= 108'o2737_4551_0202_4374_0007_0700_0000_0077_7740;
            12'o1025: crom <= 108'o2715_3443_0300_4174_4007_0700_0200_0003_0012;
            12'o1026: crom <= 108'o0534_4443_0000_4174_4007_0630_2000_0060_0000;
            12'o1027: crom <= 108'o2442_4553_0300_4374_4007_0331_0000_0000_0001;
            12'o1030: crom <= 108'o2122_4443_0000_4174_4007_0700_0010_0000_0000;
            12'o1031: crom <= 108'o3315_3771_0003_7274_4007_0701_0000_0000_0244;
            12'o1032: crom <= 108'o3315_3440_0404_1174_4007_0700_0400_0000_1443;
            12'o1033: crom <= 108'o1036_3444_0505_4174_4007_0700_0000_0000_0000;
            12'o1034: crom <= 108'o2716_3441_0302_4174_4617_0700_0000_0000_0100;
            12'o1035: crom <= 108'o1034_3333_0002_4174_4167_0700_0000_0000_0000;
            12'o1036: crom <= 108'o1064_3440_0505_0174_4007_0700_0400_0000_0000;
            12'o1037: crom <= 108'o0003_3441_0503_4174_4004_1700_0000_0000_0000;
            12'o1040: crom <= 108'o2642_3771_0003_7274_4007_0622_0010_0000_0423;
            12'o1041: crom <= 108'o2642_3771_0003_7274_4007_0622_0010_0000_0424;
            12'o1042: crom <= 108'o1047_3333_0004_7174_4007_0700_0400_0000_0423;
            12'o1043: crom <= 108'o1047_3333_0004_7174_4007_0700_0400_0000_0424;
            12'o1044: crom <= 108'o0220_3333_0005_4175_5003_7701_0200_0000_0002;
            12'o1045: crom <= 108'o2720_3333_0005_4175_5007_0701_0200_0000_0002;
            12'o1046: crom <= 108'o0614_3776_0005_0274_4007_0631_0000_0000_0000;
            12'o1047: crom <= 108'o1130_0113_0405_4174_4007_0700_0200_0024_1016;
            12'o1050: crom <= 108'o0560_3771_0004_1276_6007_0701_0010_0000_1444;
            12'o1051: crom <= 108'o3331_3771_0005_1276_6007_0701_0000_0000_1444;
            12'o1052: crom <= 108'o0460_4443_0000_4174_4007_0700_0000_0000_0000;
            12'o1053: crom <= 108'o0642_0113_0505_0174_4007_0521_0400_0000_0000;
            12'o1054: crom <= 108'o1264_5002_0000_4174_4007_0621_0010_0000_0000;
            12'o1055: crom <= 108'o2466_3771_0004_2274_4007_0120_0000_0000_0000;
            12'o1056: crom <= 108'o3247_3446_1200_4174_4007_0700_0000_0000_0000;
            12'o1057: crom <= 108'o0001_3771_0003_7274_4124_1701_0000_0000_0422;
            12'o1060: crom <= 108'o1060_3773_0000_4304_4003_1702_0000_0000_0000;
            12'o1061: crom <= 108'o1503_3333_0005_7174_4007_0700_0400_0000_0213;
            12'o1062: crom <= 108'o3556_4553_0500_4374_4007_0321_0010_0076_0740;
            12'o1063: crom <= 108'o3724_3771_0006_4374_4007_0700_0000_0000_0000;
            12'o1064: crom <= 108'o0100_3223_0000_1174_4156_4700_0400_0000_1441;
            12'o1065: crom <= 108'o1501_4571_1206_4374_4007_0700_0000_0037_0000;
            12'o1066: crom <= 108'o3257_4521_0206_4374_4007_0700_0000_0000_0740;
            12'o1067: crom <= 108'o1501_4571_1206_4374_4007_0700_0000_0037_0000;
            12'o1070: crom <= 108'o3727_3333_0005_7174_4007_0700_0400_0000_0213;
            12'o1071: crom <= 108'o1503_3333_0005_7174_4007_0700_0400_0000_0213;
            12'o1072: crom <= 108'o3727_3333_0005_7174_4007_0700_0400_0000_0213;
            12'o1073: crom <= 108'o3727_3333_0005_7174_4007_0700_0400_0000_0213;
            12'o1074: crom <= 108'o2274_3333_0003_7174_4007_0520_0410_0000_0242;
            12'o1075: crom <= 108'o0001_4221_0013_4170_4004_1700_0000_0000_0000;
            12'o1076: crom <= 108'o0716_4443_0000_7174_4003_7700_0000_0000_0241;
            12'o1077: crom <= 108'o0644_4443_0000_4174_4007_0630_2000_0060_0000;
            12'o1100: crom <= 108'o2702_4221_0013_4170_4007_0370_0000_0000_0000;
            12'o1101: crom <= 108'o3167_3771_0003_7274_4007_0701_0000_0000_0212;
            12'o1102: crom <= 108'o1562_0111_0701_4174_4007_0700_0000_0000_0000;
            12'o1103: crom <= 108'o3463_3771_0013_4370_4007_0700_0000_0000_0011;
            12'o1104: crom <= 108'o3463_3771_0013_4370_4007_0700_0000_0000_0012;
            12'o1105: crom <= 108'o2310_3771_0013_4370_4007_0700_0000_0000_0003;
            12'o1106: crom <= 108'o3472_3771_0013_4370_4007_0700_0000_0000_0012;
            12'o1107: crom <= 108'o3467_3771_0013_4370_4007_0700_0000_0000_0011;
            12'o1110: crom <= 108'o3461_3771_0013_4370_4007_0700_0000_0000_0011;
            12'o1111: crom <= 108'o2302_4221_0013_4170_4007_0700_0000_0000_0000;
            12'o1112: crom <= 108'o2310_4221_0013_4170_4007_0700_0000_0000_0000;
            12'o1113: crom <= 108'o2310_3771_0013_4370_4007_0700_0000_0000_0011;
            12'o1114: crom <= 108'o3661_0111_0702_4170_4007_0700_0210_0004_0012;
            12'o1115: crom <= 108'o3572_4551_0404_4370_4007_0700_0010_0077_0000;
            12'o1116: crom <= 108'o1123_4551_0303_0274_4007_0700_0000_0000_0000;
            12'o1117: crom <= 108'o1400_3333_0004_7174_4007_0700_0400_0000_0301;
            12'o1120: crom <= 108'o3561_3771_0003_7274_4117_0700_0010_0000_0301;
            12'o1121: crom <= 108'o3577_3333_0002_4174_4007_0700_0200_0003_0012;
            12'o1122: crom <= 108'o1764_4443_0000_4174_4007_0700_0000_0000_0000;
            12'o1123: crom <= 108'o0014_3440_0303_0174_4007_0700_0400_0000_0000;
            12'o1124: crom <= 108'o3657_3333_0016_7174_4127_0700_0400_0000_0210;
            12'o1125: crom <= 108'o1124_4443_0000_4174_4006_7653_2000_0060_0000;
            12'o1126: crom <= 108'o3657_3333_0016_7174_4127_0700_0400_0000_0210;
            12'o1127: crom <= 108'o2473_3333_0016_7174_4007_0700_0400_0000_0210;
            12'o1130: crom <= 108'o3767_3771_0003_4365_5007_0700_0210_0000_0002;
            12'o1131: crom <= 108'o1134_4553_0300_4374_4007_0321_0000_0000_0077;
            12'o1132: crom <= 108'o2561_0551_0303_7274_4007_0701_0000_0000_0215;
            12'o1133: crom <= 108'o2566_3770_0305_4344_4007_0670_0000_0000_0000;
            12'o1134: crom <= 108'o2672_4553_1300_4374_4007_0321_0000_0001_0000;
            12'o1135: crom <= 108'o2622_4251_0304_4374_4007_0700_0010_0000_3777;
            12'o1136: crom <= 108'o1143_4443_0000_4174_4007_0700_0200_0003_0002;
            12'o1137: crom <= 108'o3737_3551_0606_4374_0007_0700_0000_0010_0000;
            12'o1140: crom <= 108'o3561_3771_0003_7274_4117_0701_0010_0000_0301;
            12'o1141: crom <= 108'o2673_4443_0000_4174_4007_0700_0000_0000_0000;
            12'o1142: crom <= 108'o1507_4223_0000_4364_4277_0700_0200_0000_0010;
            12'o1143: crom <= 108'o1477_3333_0003_4175_5007_0701_0200_0000_0002;
            12'o1144: crom <= 108'o2724_3443_0300_4174_4007_0700_0200_0003_0312;
            12'o1145: crom <= 108'o2723_3443_0300_4174_4007_0700_0200_0003_0312;
            12'o1146: crom <= 108'o1147_4443_0000_4174_4467_0700_0000_0001_2000;
            12'o1147: crom <= 108'o0221_3771_0001_4361_5007_0700_0200_0000_0002;
            12'o1150: crom <= 108'o1152_0113_0503_0174_4407_0521_0400_0000_0000;
            12'o1151: crom <= 108'o1154_0113_0503_0174_4407_0521_0400_0000_0000;
            12'o1152: crom <= 108'o0100_4443_0000_4174_4156_4700_0000_0000_0000;
            12'o1153: crom <= 108'o0555_4443_0000_4174_4467_0700_0000_0001_2000;
            12'o1154: crom <= 108'o0555_4443_0000_4174_4467_0700_0000_0001_2000;
            12'o1155: crom <= 108'o0100_4443_0000_4174_4156_4700_0000_0000_0000;
            12'o1156: crom <= 108'o1510_0111_1104_4174_4007_0700_0010_0000_0000;
            12'o1157: crom <= 108'o1160_3333_0010_4174_4007_0520_0000_0000_0000;
            12'o1160: crom <= 108'o0310_3333_0004_4174_4007_0700_0200_0021_1016;
            12'o1161: crom <= 108'o1162_3770_0203_4344_4007_0700_0000_0000_0000;
            12'o1162: crom <= 108'o2745_4521_1203_4074_0007_0700_0010_0000_0000;
            12'o1163: crom <= 108'o0314_3333_0004_4174_4007_0700_0200_0021_1016;
            12'o1164: crom <= 108'o1165_3551_0505_4370_4007_0700_0000_0000_0001;
            12'o1165: crom <= 108'o1166_4553_0300_4374_4007_0321_0000_0001_0000;
            12'o1166: crom <= 108'o1167_3551_0505_4370_4007_0700_0000_0000_0004;
            12'o1167: crom <= 108'o2743_3333_0005_4174_4007_0700_0200_0024_1016;
            12'o1170: crom <= 108'o2753_0551_0303_0274_4467_0702_4000_0001_0001;
            12'o1171: crom <= 108'o2752_7441_1205_4174_4007_0700_0000_0000_0000;
            12'o1172: crom <= 108'o2753_2551_0303_0274_4467_0702_0000_0001_0001;
            12'o1173: crom <= 108'o2753_2551_0303_0274_4467_0702_4000_0001_0001;
            12'o1174: crom <= 108'o1404_4551_0404_4374_0007_0700_0000_0037_7777;
            12'o1175: crom <= 108'o1404_3551_0404_4374_0007_0700_0000_0040_0000;
            12'o1176: crom <= 108'o2755_3445_0404_4174_4007_0700_0000_0000_0000;
            12'o1177: crom <= 108'o1500_3221_0003_4174_4003_7700_0200_0003_0001;
            12'o1200: crom <= 108'o1202_3770_0404_4174_0007_0520_0000_0000_0000;
            12'o1201: crom <= 108'o1500_7001_0003_4174_4003_7700_0200_0003_0001;
            12'o1202: crom <= 108'o1404_3221_0003_4174_4467_0700_0000_0041_1000;
            12'o1203: crom <= 108'o1404_7001_0003_4174_4467_0700_0000_0041_1000;
            12'o1204: crom <= 108'o1500_4001_0004_4174_4003_7700_0200_0003_0001;
            12'o1205: crom <= 108'o1206_4113_0616_4174_4007_0520_0000_0000_0000;
            12'o1206: crom <= 108'o1500_7001_0004_4174_4003_7700_0200_0003_0001;
            12'o1207: crom <= 108'o1404_7001_0004_4174_4467_0700_0000_0041_1000;
            12'o1210: crom <= 108'o2773_3223_0000_1174_4007_0700_0400_0000_1441;
            12'o1211: crom <= 108'o2767_7003_0000_1174_4007_0700_0400_0000_1441;
            12'o1212: crom <= 108'o0110_3443_0100_4174_4156_4700_0200_0014_0012;
            12'o1213: crom <= 108'o1400_4443_0000_4174_4467_0700_0000_0041_1000;
            12'o1214: crom <= 108'o0161_4221_0003_4174_4007_0700_0000_0000_0000;
            12'o1215: crom <= 108'o0161_2441_0703_4174_4007_0700_4000_0000_0000;
            12'o1216: crom <= 108'o3007_3441_0306_4174_4007_0700_0000_0000_0000;
            12'o1217: crom <= 108'o0164_3333_0005_4174_4007_0621_0000_0000_0000;
            12'o1220: crom <= 108'o1222_2113_0305_4174_4007_0521_4000_0000_0000;
            12'o1221: crom <= 108'o1222_0113_0305_4174_4007_0521_0000_0000_0000;
            12'o1222: crom <= 108'o0555_4443_0000_4174_4467_0700_0000_0051_1000;
            12'o1223: crom <= 108'o0161_3441_0603_4174_4007_0700_0000_0000_0000;
            12'o1224: crom <= 108'o1230_3446_0505_4174_4007_0700_0000_0000_0000;
            12'o1225: crom <= 108'o1226_3446_0505_4174_4007_0520_0000_0000_0000;
            12'o1226: crom <= 108'o1230_4003_0000_4174_4007_0621_0000_0000_0000;
            12'o1227: crom <= 108'o3012_4751_1217_4374_4007_0700_0000_0000_0005;
            12'o1230: crom <= 108'o3015_3446_0505_4174_4047_0700_0000_0000_0000;
            12'o1231: crom <= 108'o0555_4443_0000_4174_4467_0700_0000_0051_1000;
            12'o1232: crom <= 108'o3042_3446_0303_4174_4007_0700_0010_0000_0000;
            12'o1233: crom <= 108'o1234_2113_0305_4174_4007_0521_4000_0000_0000;
            12'o1234: crom <= 108'o1236_2113_0305_4174_4007_0620_4000_0000_0000;
            12'o1235: crom <= 108'o3020_3221_0004_4174_4007_0700_0000_0000_0000;
            12'o1236: crom <= 108'o0033_3333_0017_4174_4003_5701_0000_0000_0000;
            12'o1237: crom <= 108'o1240_1003_0600_4174_4007_0521_4000_0000_0000;
            12'o1240: crom <= 108'o0033_3333_0017_4174_4003_5701_0000_0000_0000;
            12'o1241: crom <= 108'o3020_3221_0004_4174_4007_0700_0000_0000_0000;
            12'o1242: crom <= 108'o3042_3442_0400_4174_4007_0700_0010_0000_0000;
            12'o1243: crom <= 108'o3023_3221_0004_4174_4007_0700_0000_0000_0000;
            12'o1244: crom <= 108'o3030_3440_1616_1174_4007_0700_0400_0000_1441;
            12'o1245: crom <= 108'o3032_4223_0000_1174_4007_0700_0400_0000_1441;
            12'o1246: crom <= 108'o3036_3442_0400_4174_4007_0700_0000_0000_0000;
            12'o1247: crom <= 108'o3033_0112_0406_4174_4007_0700_0000_0000_0000;
            12'o1250: crom <= 108'o0100_4003_0000_1174_4156_4700_0400_0000_1443;
            12'o1251: crom <= 108'o3041_4002_0000_1174_4007_0700_0000_0000_1443;
            12'o1252: crom <= 108'o3045_4221_0004_4174_4007_0700_0000_0000_0000;
            12'o1253: crom <= 108'o1254_2222_0000_4174_4007_0621_4000_0000_0000;
            12'o1254: crom <= 108'o3044_7441_0303_4174_4007_0700_0000_0000_0000;
            12'o1255: crom <= 108'o3044_2441_0303_4174_4007_0700_4000_0000_0000;
            12'o1256: crom <= 108'o3047_3446_0303_4174_4007_0700_0000_0000_0000;
            12'o1257: crom <= 108'o3046_2441_0505_4174_4007_0700_4000_0000_0000;
            12'o1260: crom <= 108'o1260_0114_0503_4174_4067_0630_2100_0060_0000;
            12'o1261: crom <= 108'o3053_3444_1717_4174_4067_0700_0100_0000_0000;
            12'o1262: crom <= 108'o3054_3444_0303_4174_4007_0700_0000_0000_0000;
            12'o1263: crom <= 108'o1262_0111_0503_4174_4007_0700_0000_0000_0000;
            12'o1264: crom <= 108'o3057_1114_0604_4174_4057_0700_4000_0000_0000;
            12'o1265: crom <= 108'o3057_0114_0604_4174_4057_0700_0000_0000_0000;
            12'o1266: crom <= 108'o3057_0114_0604_4174_4067_0700_0100_0000_0000;
            12'o1267: crom <= 108'o0002_4444_0002_4174_4064_1700_0100_0000_0000;
            12'o1270: crom <= 108'o3064_7772_0000_1274_4007_0701_0000_0000_1442;
            12'o1271: crom <= 108'o3062_1772_0000_1274_4007_0701_4000_0000_1442;
            12'o1272: crom <= 108'o3065_7772_0000_1274_4007_0701_0000_0000_1441;
            12'o1273: crom <= 108'o3063_1772_0000_1274_4007_0701_4000_0000_1441;
            12'o1274: crom <= 108'o3066_7771_0003_0274_4007_0700_0000_0000_0000;
            12'o1275: crom <= 108'o3066_1771_0003_0274_4007_0701_4000_0000_0000;
            12'o1276: crom <= 108'o2220_7441_0303_4174_4467_0700_0000_0001_0001;
            12'o1277: crom <= 108'o2220_2441_0303_4174_4467_0701_4000_0001_0001;
            12'o1300: crom <= 108'o2220_7441_0303_4174_4007_0700_0000_0000_0000;
            12'o1301: crom <= 108'o2220_2441_0303_4174_4007_0700_4000_0000_0000;
            12'o1302: crom <= 108'o1302_3447_0404_4174_4007_0630_2000_0060_0000;
            12'o1303: crom <= 108'o3130_4557_0404_4374_4007_0701_0000_0000_0176;
            12'o1304: crom <= 108'o1304_3447_0505_4174_4007_0630_2000_0060_0000;
            12'o1305: crom <= 108'o1306_3333_0005_7174_4007_0621_0400_0000_0222;
            12'o1306: crom <= 108'o0660_3442_0400_4174_4007_0700_2000_0071_0042;
            12'o1307: crom <= 108'o1404_3771_0003_7274_4007_0701_0000_0000_0223;
            12'o1310: crom <= 108'o0570_0662_0000_0274_4007_0522_2000_0071_0042;
            12'o1311: crom <= 108'o0555_4443_0000_4174_4467_0700_0000_0051_1000;
            12'o1312: crom <= 108'o3145_0661_0005_7274_4407_0701_0000_0000_0223;
            12'o1313: crom <= 108'o3144_1002_0700_4170_4007_0700_4000_0000_0000;
            12'o1314: crom <= 108'o1314_3445_0303_4174_4007_0630_2000_0060_0000;
            12'o1315: crom <= 108'o3152_4551_0505_4374_0007_0700_0000_0000_7777;
            12'o1316: crom <= 108'o3663_3443_0400_4174_4007_0700_0210_0004_0712;
            12'o1317: crom <= 108'o3154_4221_0006_4174_0007_0700_0000_0000_0000;
            12'o1320: crom <= 108'o3164_3443_0600_4174_4007_0700_0200_0003_0312;
            12'o1321: crom <= 108'o3162_3443_0600_4174_4007_0700_0200_0003_0312;
            12'o1322: crom <= 108'o3165_4443_0000_4174_4007_0700_0000_0000_0000;
            12'o1323: crom <= 108'o1324_2113_0603_4174_4007_0521_4000_0000_0000;
            12'o1324: crom <= 108'o1400_4221_0013_4170_4007_0700_0000_0000_0000;
            12'o1325: crom <= 108'o1326_0111_0704_4174_4007_0370_0000_0000_0000;
            12'o1326: crom <= 108'o3162_0111_0706_4170_4007_0700_0200_0003_0312;
            12'o1327: crom <= 108'o3164_0111_0706_4170_4007_0700_0200_0003_0312;
            12'o1330: crom <= 108'o1400_4221_0013_4170_4007_0700_0000_0000_0000;
            12'o1331: crom <= 108'o3166_0111_0706_4174_4007_0700_0000_0000_0000;
            12'o1332: crom <= 108'o3175_4551_0303_4374_0007_0700_0000_0000_0777;
            12'o1333: crom <= 108'o3175_3551_0303_4374_0007_0700_0000_0077_7000;
            12'o1334: crom <= 108'o3175_4551_0505_4374_0007_0700_0000_0000_0777;
            12'o1335: crom <= 108'o3175_3551_0505_4374_0007_0700_0000_0077_7000;
            12'o1336: crom <= 108'o1336_3446_0505_4174_4047_0630_2000_0060_0000;
            12'o1337: crom <= 108'o0420_0111_0503_4174_4003_4701_0000_0000_0000;
            12'o1340: crom <= 108'o3176_4551_0606_4374_0007_0700_0000_0000_0777;
            12'o1341: crom <= 108'o3176_3551_0606_4374_0007_0700_0000_0077_7000;
            12'o1342: crom <= 108'o1344_3771_0003_0276_6007_0520_1000_0030_2000;
            12'o1343: crom <= 108'o0555_4443_0000_4174_4467_0700_0000_0071_1000;
            12'o1344: crom <= 108'o3201_4551_0303_4374_0007_0700_0000_0000_0777;
            12'o1345: crom <= 108'o3202_3551_0303_4374_0007_0700_0000_0077_7000;
            12'o1346: crom <= 108'o1350_2113_0406_4174_4007_0311_4000_0000_0000;
            12'o1347: crom <= 108'o1346_2445_0506_4174_4007_0700_4000_0000_0000;
            12'o1350: crom <= 108'o1352_3447_0606_4174_4007_0700_0000_0000_0000;
            12'o1351: crom <= 108'o0555_4443_0000_4174_4467_0700_0000_0071_1000;
            12'o1352: crom <= 108'o3665_3445_0303_4174_4007_0700_0010_0000_0000;
            12'o1353: crom <= 108'o0144_2113_0604_4174_4007_0421_4000_0000_0000;
            12'o1354: crom <= 108'o1356_2441_0305_4174_4007_0521_4000_0000_0000;
            12'o1355: crom <= 108'o1363_4222_0000_4174_4007_0700_1000_0071_0233;
            12'o1356: crom <= 108'o1360_4553_0500_4374_4007_0321_0000_0077_7000;
            12'o1357: crom <= 108'o3205_4222_0000_4174_4007_0700_1000_0071_0244;
            12'o1360: crom <= 108'o3205_4222_0000_4174_4007_0700_1000_0071_0244;
            12'o1361: crom <= 108'o1363_4222_0000_4174_4007_0700_1000_0071_0233;
            12'o1362: crom <= 108'o1362_3446_0303_4174_4047_0630_2000_0060_0000;
            12'o1363: crom <= 108'o0420_3333_0003_4174_4003_4701_0000_0000_0000;
            12'o1364: crom <= 108'o1363_4551_0303_4374_0007_0700_0000_0000_0777;
            12'o1365: crom <= 108'o1363_3551_0303_4374_0007_0700_0000_0077_7000;
            12'o1366: crom <= 108'o1366_3446_0303_4174_4047_0630_2000_0060_0000;
            12'o1367: crom <= 108'o0063_3447_0705_4174_4003_7700_0000_0000_0000;
            12'o1370: crom <= 108'o1370_3445_0303_4174_4007_0630_2000_0060_0000;
            12'o1371: crom <= 108'o0100_3440_0303_0174_4156_4700_0400_0000_0000;
            12'o1372: crom <= 108'o0100_3440_0303_0174_4156_4700_0400_0000_0000;
            12'o1373: crom <= 108'o1374_3223_0000_4174_4007_0621_0000_0000_0000;
            12'o1374: crom <= 108'o1514_0111_0703_4174_4003_7700_0200_0003_0001;
            12'o1375: crom <= 108'o0073_7441_1205_4174_4007_0700_0000_0000_0000;
            12'o1376: crom <= 108'o0420_3444_0303_4174_4063_4701_1000_0041_1777;
            12'o1377: crom <= 108'o1514_4443_0000_4174_4003_7700_0200_0003_0001;
            12'o1400: crom <= 108'o0110_3443_0100_4174_4156_4700_0200_0014_0012;
            12'o1401: crom <= 108'o0110_0111_0701_4170_4156_4700_0200_0014_0012;
            12'o1402: crom <= 108'o1500_3770_0303_4344_4003_7700_0200_0003_0001;
            12'o1403: crom <= 108'o1404_3333_0003_4174_4007_0520_0000_0000_0000;
            12'o1404: crom <= 108'o1500_4443_0000_4174_4003_7700_0200_0003_0001;
            12'o1405: crom <= 108'o1404_2441_0303_4174_4467_0701_4000_0001_0001;
            12'o1406: crom <= 108'o0506_3771_0005_0276_6007_0700_0200_0003_0002;
            12'o1407: crom <= 108'o1500_3771_0003_0276_0003_7700_0200_0003_0001;
            12'o1410: crom <= 108'o1500_3771_0003_0270_6003_7700_0200_0003_0001;
            12'o1411: crom <= 108'o1410_3770_0303_4344_4007_0700_0000_0000_0000;
            12'o1412: crom <= 108'o1407_3770_0303_4344_4007_0700_0000_0000_0000;
            12'o1413: crom <= 108'o0511_3770_0303_4344_4007_0700_0000_0000_0000;
            12'o1414: crom <= 108'o1500_3770_0303_4344_0003_7700_0200_0003_0001;
            12'o1415: crom <= 108'o0512_3770_0303_4344_4007_0700_0000_0000_0000;
            12'o1416: crom <= 108'o1500_3770_0303_4340_4003_7700_0200_0003_0001;
            12'o1417: crom <= 108'o1420_3333_0003_4174_4007_0530_0000_0000_0000;
            12'o1420: crom <= 108'o1500_5731_0003_4174_4003_7700_0200_0003_0001;
            12'o1421: crom <= 108'o1500_5431_1203_4174_4003_7700_0200_0003_0001;
            12'o1422: crom <= 108'o1424_3333_0003_4174_4007_0530_0000_0000_0000;
            12'o1423: crom <= 108'o1426_3333_0003_4174_4007_0520_0000_0000_0000;
            12'o1424: crom <= 108'o1402_3771_0003_4374_0007_0700_0000_0000_0000;
            12'o1425: crom <= 108'o1402_3771_0003_4374_0007_0700_0000_0077_7777;
            12'o1426: crom <= 108'o1402_3771_0003_4370_4007_0700_0000_0000_0000;
            12'o1427: crom <= 108'o1402_3771_0003_4370_4007_0700_0000_0077_7777;
            12'o1430: crom <= 108'o1432_3333_0003_4174_4007_0520_0000_0000_0000;
            12'o1431: crom <= 108'o1136_0111_0703_4174_4467_0701_0000_0001_0001;
            12'o1432: crom <= 108'o1500_5371_0003_4174_4003_7700_0200_0003_0001;
            12'o1433: crom <= 108'o1500_5341_1203_4174_4003_7700_0200_0003_0001;
            12'o1434: crom <= 108'o3070_4551_0404_4374_0007_0700_0010_0037_7777;
            12'o1435: crom <= 108'o2660_4553_0400_4374_4007_0331_0000_0002_0000;
            12'o1436: crom <= 108'o1515_3440_0404_1174_4007_0700_0400_0000_1441;
            12'o1437: crom <= 108'o1136_1111_0703_4174_4467_0701_4000_0001_0001;
            12'o1440: crom <= 108'o0270_3771_0005_0276_6003_7700_0000_0000_0000;
            12'o1441: crom <= 108'o1500_4221_0003_4174_4003_7700_0200_0003_0001;
            12'o1442: crom <= 108'o1500_4551_0303_0274_4003_7700_0200_0003_0001;
            12'o1443: crom <= 108'o1500_5551_0303_0274_4003_7700_0200_0003_0001;
            12'o1444: crom <= 108'o1442_7441_0303_4174_4007_0700_0000_0000_0000;
            12'o1445: crom <= 108'o1500_6551_0303_0274_4003_7700_0200_0003_0001;
            12'o1446: crom <= 108'o1500_3551_0303_0274_4003_7700_0200_0003_0001;
            12'o1447: crom <= 108'o1443_7441_0303_4174_4007_0700_0000_0000_0000;
            12'o1450: crom <= 108'o1500_7551_0303_0274_4003_7700_0200_0003_0001;
            12'o1451: crom <= 108'o1500_7771_0003_0274_4003_7700_0200_0003_0001;
            12'o1452: crom <= 108'o0564_7771_0005_0274_4007_0700_0000_0000_0000;
            12'o1453: crom <= 108'o1500_7441_0303_4174_4003_7700_0200_0003_0001;
            12'o1454: crom <= 108'o1446_7441_0303_4174_4007_0700_0000_0000_0000;
            12'o1455: crom <= 108'o1453_4551_0303_0274_4007_0700_0000_0000_0000;
            12'o1456: crom <= 108'o1500_2441_0703_4174_4003_7700_4200_0003_0001;
            12'o1457: crom <= 108'o1170_0551_0404_1274_4007_0562_0000_0000_1441;
            12'o1460: crom <= 108'o2436_4443_0000_4174_4007_0700_0010_0000_0000;
            12'o1461: crom <= 108'o2446_3771_0005_0276_6007_0700_0000_0000_0000;
            12'o1462: crom <= 108'o0502_4551_1205_0276_6007_0622_0000_0000_0000;
            12'o1463: crom <= 108'o1400_3440_0303_0174_4007_0700_0400_0000_0000;
            12'o1464: crom <= 108'o0544_4443_0000_4174_4007_0630_2000_0060_0000;
            12'o1465: crom <= 108'o1026_3333_0003_4174_4007_0700_2000_0031_5777;
            12'o1466: crom <= 108'o0554_3333_0003_4174_4007_0330_3000_0041_4000;
            12'o1467: crom <= 108'o1062_3771_0005_4365_5007_0700_0200_0000_0002;
            12'o1470: crom <= 108'o0742_4443_0000_4174_4007_0630_2000_0060_0000;
            12'o1471: crom <= 108'o1077_3333_0003_4174_4007_0700_2000_0031_5777;
            12'o1472: crom <= 108'o1473_3770_0303_4344_4007_0700_0000_0000_0000;
            12'o1473: crom <= 108'o0014_4221_0005_4174_4003_7700_0000_0000_0000;
            12'o1474: crom <= 108'o1475_3770_0303_4344_4007_0700_0000_0000_0000;
            12'o1475: crom <= 108'o0014_4551_0305_0274_4003_7700_0000_0000_0000;
            12'o1476: crom <= 108'o0250_2551_0303_0274_4003_7701_4000_0000_0000;
            12'o1477: crom <= 108'o0744_3770_0303_4174_0007_0360_0000_0000_0000;
            12'o1500: crom <= 108'o2607_3551_0606_4374_4007_0700_0000_0004_0000;
            12'o1501: crom <= 108'o2670_3333_0005_7174_4007_0700_0400_0000_0213;
            12'o1502: crom <= 108'o2656_3111_0506_4174_4007_0700_0000_0000_0000;
            12'o1503: crom <= 108'o1140_4443_0000_4174_4007_0370_0000_0000_0000;
            12'o1504: crom <= 108'o0434_4443_0000_4174_4007_0360_0000_0000_0000;
            12'o1505: crom <= 108'o1515_3440_0404_1174_4007_0700_0400_0000_1441;
            12'o1506: crom <= 108'o1505_3333_0003_4175_5007_0701_0200_0000_0002;
            12'o1507: crom <= 108'o3762_3771_0003_7274_4007_0701_0000_0000_0210;
            12'o1510: crom <= 108'o0001_4223_0000_4364_4274_1700_0200_0000_0010;
            12'o1511: crom <= 108'o2700_3333_0003_4174_4467_0700_0000_0000_0004;
            12'o1512: crom <= 108'o2704_3443_0300_4174_4007_0700_0200_0021_1016;
            12'o1513: crom <= 108'o1563_3333_0005_4175_5007_0701_0200_0000_0002;
            12'o1514: crom <= 108'o0104_4751_1217_4374_4007_0700_0000_0000_1000;
            12'o1515: crom <= 108'o0100_3440_0303_0174_4156_4700_0400_0000_0000;
            12'o1516: crom <= 108'o1400_3333_0003_4175_5007_0701_0200_0000_0002;
            12'o1517: crom <= 108'o1515_3333_0003_4175_5007_0701_0200_0000_0002;
            12'o1520: crom <= 108'o0110_3441_0301_4170_4156_4700_0200_0014_0012;
            12'o1521: crom <= 108'o0110_3441_0301_4170_4156_4700_0200_0014_0012;
            12'o1522: crom <= 108'o0150_1113_0701_4170_4007_0700_4200_0004_0012;
            12'o1523: crom <= 108'o2737_4551_0202_4374_0007_0700_0000_0077_7740;
            12'o1524: crom <= 108'o1004_4443_0000_4174_4007_0340_0000_0000_0000;
            12'o1525: crom <= 108'o2606_3443_0300_4174_4007_0700_0200_0004_0012;
            12'o1526: crom <= 108'o0320_4443_0000_4174_4007_0340_0000_0000_0000;
            12'o1527: crom <= 108'o1014_4443_0000_4174_4007_0340_0000_0000_0000;
            12'o1530: crom <= 108'o1010_1113_0701_4170_4007_0040_4200_0004_0012;
            12'o1531: crom <= 108'o2737_4551_0202_4374_0007_0700_0000_0077_7740;
            12'o1532: crom <= 108'o0300_1113_0701_4170_4007_0040_4200_0004_0012;
            12'o1533: crom <= 108'o2737_4551_0202_4374_0007_0700_0000_0077_7740;
            12'o1534: crom <= 108'o1024_4443_0000_4174_4007_0340_0000_0000_0000;
            12'o1535: crom <= 108'o2737_4551_0202_4374_0007_0700_0000_0077_7740;
            12'o1536: crom <= 108'o2737_4551_0202_4374_0007_0700_0000_0077_7740;
            12'o1537: crom <= 108'o2737_4551_0202_4374_0007_0700_0000_0077_7740;
            12'o1540: crom <= 108'o0762_4443_0000_4174_4467_0551_0000_0001_0010;
            12'o1541: crom <= 108'o1034_4443_0000_4174_4007_0340_0000_0000_0000;
            12'o1542: crom <= 108'o0270_2551_0705_0274_4463_7702_4000_0001_0001;
            12'o1543: crom <= 108'o2717_3771_0005_4365_5007_0700_0200_0000_0002;
            12'o1544: crom <= 108'o2717_3741_0105_4074_4467_0700_0000_0005_0000;
            12'o1545: crom <= 108'o2721_3771_0004_0276_6007_0701_0200_0004_0712;
            12'o1546: crom <= 108'o2725_3771_0004_0276_6007_0701_0200_0004_0712;
            12'o1547: crom <= 108'o0270_0551_1505_0274_4403_7701_0000_0000_0000;
            12'o1550: crom <= 108'o2727_3741_0105_4074_4007_0700_0000_0000_0000;
            12'o1551: crom <= 108'o2726_3770_0303_4344_0007_0700_0000_0000_0000;
            12'o1552: crom <= 108'o2730_3741_0105_4074_4467_0700_0000_0005_0000;
            12'o1553: crom <= 108'o3713_3551_0303_4374_0007_0700_0000_0016_0000;
            12'o1554: crom <= 108'o2733_3441_0305_4174_4007_0700_0200_0003_0002;
            12'o1555: crom <= 108'o2734_3771_0005_0276_6007_0700_0000_0000_0000;
            12'o1556: crom <= 108'o2737_4551_0202_4374_0007_0700_0000_0077_7740;
            12'o1557: crom <= 108'o0400_4751_1203_4374_4007_0700_0000_0000_0040;
            12'o1560: crom <= 108'o1500_0551_0303_0274_4463_7701_0200_0001_0001;
            12'o1561: crom <= 108'o1500_2551_0303_0274_4463_7701_4200_0001_0001;
            12'o1562: crom <= 108'o2710_4221_0013_4170_4007_0370_0000_0000_0000;
            12'o1563: crom <= 108'o2743_0111_0703_4174_4007_0700_0200_0024_1016;
            12'o1564: crom <= 108'o0001_0111_0703_4170_4004_1700_0200_0023_1016;
            12'o1565: crom <= 108'o3067_3771_0004_1276_6007_0701_0010_0000_1441;
            12'o1566: crom <= 108'o2761_3447_0303_4174_4007_0700_0000_0000_0000;
            12'o1567: crom <= 108'o0531_0113_0207_4174_4007_0700_0200_0003_0312;
            12'o1570: crom <= 108'o1340_3771_0006_0276_6007_0521_1000_0040_2000;
            12'o1571: crom <= 108'o2756_3442_0300_0174_4007_0700_0000_0000_0000;
            12'o1572: crom <= 108'o0000_0000_0000_0000_0000_0000_0000_0000_0000;
            12'o1573: crom <= 108'o0000_0000_0000_0000_0000_0000_0000_0000_0000;
            12'o1574: crom <= 108'o1342_3441_0305_0174_4007_0621_0000_0000_0000;
            12'o1575: crom <= 108'o0000_0000_0000_0000_0000_0000_0000_0000_0000;
            12'o1576: crom <= 108'o1577_2441_0303_4174_4007_0700_4000_0000_0000;
            12'o1577: crom <= 108'o0670_3771_0005_0276_6006_7701_2000_0020_2000;
            12'o1600: crom <= 108'o3003_3441_0305_0174_4007_0700_0000_0000_0000;
            12'o1601: crom <= 108'o3004_3441_0305_4174_4007_0700_0000_0000_0000;
            12'o1602: crom <= 108'o0000_0000_0000_0000_0000_0000_0000_0000_0000;
            12'o1603: crom <= 108'o0000_0000_0000_0000_0000_0000_0000_0000_0000;
            12'o1604: crom <= 108'o0000_0000_0000_0000_0000_0000_0000_0000_0000;
            12'o1605: crom <= 108'o0000_0000_0000_0000_0000_0000_0000_0000_0000;
            12'o1606: crom <= 108'o0000_0000_0000_0000_0000_0000_0000_0000_0000;
            12'o1607: crom <= 108'o0000_0000_0000_0000_0000_0000_0000_0000_0000;
            12'o1610: crom <= 108'o0240_4443_0000_4174_4007_0360_0000_0000_0000;
            12'o1611: crom <= 108'o0270_0551_0705_0274_4463_7702_0000_0001_0001;
            12'o1612: crom <= 108'o0572_3771_0003_0276_6007_0700_1000_0031_1777;
            12'o1613: crom <= 108'o0611_4551_1203_0276_6007_0700_1000_0041_0001;
            12'o1614: crom <= 108'o2436_4443_0000_4174_4007_0700_0010_0000_0000;
            12'o1615: crom <= 108'o1172_2551_0404_1274_4007_0562_4000_0000_1441;
            12'o1616: crom <= 108'o1354_4553_0300_4374_4007_0321_0000_0077_7000;
            12'o1617: crom <= 108'o0014_4551_0305_0274_4003_7700_0000_0000_0000;
            12'o1620: crom <= 108'o0350_3770_0305_4334_4016_7351_0010_0033_6000;
            12'o1621: crom <= 108'o3206_3333_0003_4174_4007_0700_2000_0041_4000;
            12'o1622: crom <= 108'o0632_4222_0000_4174_4007_0700_0000_0000_0000;
            12'o1623: crom <= 108'o0611_3771_0003_0276_6007_0700_1000_0041_0001;
            12'o1624: crom <= 108'o3077_3333_0003_4174_4217_0701_1010_0073_0500;
            12'o1625: crom <= 108'o0604_3443_0100_4174_4007_0700_0200_0014_0012;
            12'o1626: crom <= 108'o0674_4222_0000_4174_4006_7701_0000_0041_1534;
            12'o1627: crom <= 108'o3011_4112_0400_4174_4007_0700_0000_0000_0000;
            12'o1630: crom <= 108'o0350_3770_0305_4334_4016_7351_0010_0033_6000;
            12'o1631: crom <= 108'o2020_3442_0400_4174_4007_0700_2000_0071_0006;
            12'o1632: crom <= 108'o0747_3777_0003_0274_4007_0701_1000_0031_1777;
            12'o1633: crom <= 108'o0646_3777_0003_0274_4007_0701_1000_0041_0001;
            12'o1634: crom <= 108'o3072_3775_0004_0274_4007_0701_0000_0000_0000;
            12'o1635: crom <= 108'o3212_2441_0404_4174_4007_0700_4000_0000_0000;
            12'o1636: crom <= 108'o0132_3441_0406_4174_4007_0700_0000_0000_0000;
            12'o1637: crom <= 108'o3213_4557_0006_1274_4007_0701_0000_0000_1441;
            12'o1640: crom <= 108'o3153_3771_0006_0276_6007_0700_0010_0000_0000;
            12'o1641: crom <= 108'o2754_3441_0306_0174_4007_0700_0000_0000_0000;
            12'o1642: crom <= 108'o3662_3440_0505_0174_4007_0700_0410_0000_0000;
            12'o1643: crom <= 108'o3161_0551_0405_4370_4007_0701_0000_0000_0001;
            12'o1644: crom <= 108'o2436_3441_0306_4174_4007_0700_0010_0000_0000;
            12'o1645: crom <= 108'o0000_0000_0000_0000_0000_0000_0000_0000_0000;
            12'o1646: crom <= 108'o0000_0000_0000_0000_0000_0000_0000_0000_0000;
                12'o1647: crom <= 108'o1013_3441_0305_4174_4003_7700_0000_0000_0000;
            12'o1650: crom <= 108'o2737_4551_0202_4374_0007_0700_0000_0077_7740;
            12'o1651: crom <= 108'o2737_4551_0202_4374_0007_0700_0000_0077_7740;
            12'o1652: crom <= 108'o2737_4551_0202_4374_0007_0700_0000_0077_7740;
            12'o1653: crom <= 108'o2737_4551_0202_4374_0007_0700_0000_0077_7740;
            12'o1654: crom <= 108'o2737_4551_0202_4374_0007_0700_0000_0077_7740;
            12'o1655: crom <= 108'o2737_4551_0202_4374_0007_0700_0000_0077_7740;
            12'o1656: crom <= 108'o2737_4551_0202_4374_0007_0700_0000_0077_7740;
            12'o1657: crom <= 108'o2737_4551_0202_4374_0007_0700_0000_0077_7740;
            12'o1660: crom <= 108'o2737_4551_0202_4374_0007_0700_0000_0077_7740;
            12'o1661: crom <= 108'o2737_4551_0202_4374_0007_0700_0000_0077_7740;
            12'o1662: crom <= 108'o2737_4551_0202_4374_0007_0700_0000_0077_7740;
            12'o1663: crom <= 108'o2737_4551_0202_4374_0007_0700_0000_0077_7740;
            12'o1664: crom <= 108'o2737_4551_0202_4374_0007_0700_0000_0077_7740;
            12'o1665: crom <= 108'o2737_4551_0202_4374_0007_0700_0000_0077_7740;
            12'o1666: crom <= 108'o2737_4551_0202_4374_0007_0700_0000_0077_7740;
            12'o1667: crom <= 108'o2737_4551_0202_4374_0007_0700_0000_0077_7740;
            12'o1670: crom <= 108'o0000_0000_0000_0000_0000_0000_0000_0000_0000;
            12'o1671: crom <= 108'o0000_0000_0000_0000_0000_0000_0000_0000_0000;
            12'o1672: crom <= 108'o0000_0000_0000_0000_0000_0000_0000_0000_0000;
            12'o1673: crom <= 108'o0000_0000_0000_0000_0000_0000_0000_0000_0000;
            12'o1674: crom <= 108'o0000_0000_0000_0000_0000_0000_0000_0000_0000;
            12'o1675: crom <= 108'o0000_0000_0000_0000_0000_0000_0000_0000_0000;
            12'o1676: crom <= 108'o0000_0000_0000_0000_0000_0000_0000_0000_0000;
            12'o1677: crom <= 108'o0000_0000_0000_0000_0000_0000_0000_0000_0000;
            12'o1700: crom <= 108'o0137_3771_0005_4374_4007_0700_0000_0001_0001;
            12'o1701: crom <= 108'o2737_4551_0202_4374_0007_0700_0000_0077_7740;
            12'o1702: crom <= 108'o2737_4551_0202_4374_0007_0700_0000_0077_7740;
            12'o1703: crom <= 108'o2737_4551_0202_4374_0007_0700_0000_0077_7740;
            12'o1704: crom <= 108'o3503_3771_0005_7274_4007_0701_0000_0000_0230;
            12'o1705: crom <= 108'o3516_3771_0005_7274_4007_0701_0000_0000_0230;
            12'o1706: crom <= 108'o3502_3771_0005_4304_4007_0701_0000_0000_0000;
            12'o1707: crom <= 108'o3500_3771_0005_4304_4007_0701_0000_0000_0000;
            12'o1710: crom <= 108'o2737_4551_0202_4374_0007_0700_0000_0077_7740;
            12'o1711: crom <= 108'o2737_4551_0202_4374_0007_0700_0000_0077_7740;
            12'o1712: crom <= 108'o2737_4551_0202_4374_0007_0700_0000_0077_7740;
            12'o1713: crom <= 108'o2737_4551_0202_4374_0007_0700_0000_0077_7740;
            12'o1714: crom <= 108'o2364_4553_0300_4374_4007_0331_0000_0001_0000;
            12'o1715: crom <= 108'o3613_3441_1405_4174_4007_0700_0000_0000_0000;
            12'o1716: crom <= 108'o0136_3441_1405_4174_4007_0700_0000_0000_0000;
            12'o1717: crom <= 108'o3501_3441_1405_4174_4007_0700_0000_0000_0000;
            12'o1720: crom <= 108'o2737_4551_0202_4374_0007_0700_0000_0077_7740;
            12'o1721: crom <= 108'o2352_4551_1105_4374_0007_0700_0000_0050_7700;
            12'o1722: crom <= 108'o3615_3443_0300_4174_4147_0700_0200_0000_0010;
            12'o1723: crom <= 108'o3524_3443_0300_4174_4007_0700_0200_0004_0012;
            12'o1724: crom <= 108'o2342_3445_0303_4174_4007_0700_2000_0071_0006;
            12'o1725: crom <= 108'o2350_3447_1005_4174_4007_0700_2000_0071_0006;
            12'o1726: crom <= 108'o2737_4551_0202_4374_0007_0700_0000_0077_7740;
            12'o1727: crom <= 108'o2737_4551_0202_4374_0007_0700_0000_0077_7740;
            12'o1730: crom <= 108'o2737_4551_0202_4374_0007_0700_0000_0077_7740;
            12'o1731: crom <= 108'o2737_4551_0202_4374_0007_0700_0000_0077_7740;
            12'o1732: crom <= 108'o2737_4551_0202_4374_0007_0700_0000_0077_7740;
            12'o1733: crom <= 108'o2737_4551_0202_4374_0007_0700_0000_0077_7740;
            12'o1734: crom <= 108'o2737_4551_0202_4374_0007_0700_0000_0077_7740;
            12'o1735: crom <= 108'o2737_4551_0202_4374_0007_0700_0000_0077_7740;
            12'o1736: crom <= 108'o2737_4551_0202_4374_0007_0700_0000_0077_7740;
            12'o1737: crom <= 108'o2737_4551_0202_4374_0007_0700_0000_0077_7740;
            12'o1740: crom <= 108'o0400_4751_1203_4374_4007_0700_0000_0000_0040;
            12'o1741: crom <= 108'o0400_4751_1203_4374_4007_0700_0000_0000_0040;
            12'o1742: crom <= 108'o0400_4751_1203_4374_4007_0700_0000_0000_0040;
            12'o1743: crom <= 108'o0400_4751_1203_4374_4007_0700_0000_0000_0040;
            12'o1744: crom <= 108'o0400_4751_1203_4374_4007_0700_0000_0000_0040;
            12'o1745: crom <= 108'o0000_0000_0000_0000_0000_0000_0000_0000_0000;
            12'o1746: crom <= 108'o0400_4751_1203_4374_4007_0700_0000_0000_0040;
            12'o1747: crom <= 108'o0400_4751_1203_4374_4007_0700_0000_0000_0040;
            12'o1750: crom <= 108'o0400_4751_1203_4374_4007_0700_0000_0000_0040;
            12'o1751: crom <= 108'o0400_4751_1203_4374_4007_0700_0000_0000_0040;
            12'o1752: crom <= 108'o0000_0000_0000_0000_0000_0000_0000_0000_0000;
            12'o1753: crom <= 108'o0000_0000_0000_0000_0000_0000_0000_0000_0000;
            12'o1754: crom <= 108'o3672_3443_0300_4174_4207_0700_0200_0004_0012;
            12'o1755: crom <= 108'o3673_3443_0300_4174_4207_0700_0200_0003_0012;
            12'o1756: crom <= 108'o0000_0000_0000_0000_0000_0000_0000_0000_0000;
            12'o1757: crom <= 108'o0000_0000_0000_0000_0000_0000_0000_0000_0000;
            12'o1760: crom <= 108'o3613_3771_0005_7274_4007_0701_0000_0000_0215;
            12'o1761: crom <= 108'o3613_3771_0005_7274_4007_0701_0000_0000_0216;
            12'o1762: crom <= 108'o3613_3771_0005_7274_4007_0701_0000_0000_0220;
            12'o1763: crom <= 108'o3613_3771_0005_7274_4007_0701_0000_0000_0217;
            12'o1764: crom <= 108'o3573_4451_1205_4324_4007_0700_0000_0000_0000;
            12'o1765: crom <= 108'o3613_3771_0005_7274_4007_0701_0000_0000_0302;
            12'o1766: crom <= 108'o3613_3771_0005_7274_4007_0701_0000_0000_0227;
            12'o1767: crom <= 108'o2737_4551_0202_4374_0007_0700_0000_0077_7740;
            12'o1770: crom <= 108'o3544_4443_0000_4174_4007_0703_0200_0006_0002;
            12'o1771: crom <= 108'o3546_4443_0000_4174_4007_0703_0200_0006_0002;
            12'o1772: crom <= 108'o3550_4443_0000_4174_4007_0703_0200_0006_0002;
            12'o1773: crom <= 108'o3552_4443_0000_4174_4007_0703_0200_0006_0002;
            12'o1774: crom <= 108'o3571_4443_0000_4174_4007_0700_0200_0004_0002;
            12'o1775: crom <= 108'o3602_4443_0000_4174_4007_0700_0200_0004_0002;
            12'o1776: crom <= 108'o3554_4443_0000_4174_4007_0703_0200_0006_0002;
            12'o1777: crom <= 108'o2737_4551_0202_4374_0007_0700_0000_0077_7740;
            12'o2000: crom <= 108'o0440_7441_0303_4174_4003_4701_0000_0000_0000;
            12'o2001: crom <= 108'o0440_2441_0303_4174_4003_4701_4000_0000_0000;
            12'o2002: crom <= 108'o3211_7441_0303_4174_4007_0700_0000_0000_0000;
            12'o2003: crom <= 108'o2004_3223_0000_4174_4007_0621_0000_0000_0000;
            12'o2004: crom <= 108'o3211_7441_0303_4174_4007_0700_0000_0000_0000;
            12'o2005: crom <= 108'o3211_2441_0303_4174_4007_0700_4000_0000_0000;
            12'o2006: crom <= 108'o2010_5547_0505_0374_4007_0631_0000_0077_7400;
            12'o2007: crom <= 108'o2010_3547_0505_0374_4007_0631_0000_0077_7400;
            12'o2010: crom <= 108'o2012_3442_0600_4174_4007_0700_0000_0000_0000;
            12'o2011: crom <= 108'o3215_3771_0016_0276_6007_0700_2000_0041_2000;
            12'o2012: crom <= 108'o0153_3441_0516_4174_4007_0700_0010_0000_0000;
            12'o2013: crom <= 108'o3214_3441_1605_4174_4007_0700_0000_0000_0000;
            12'o2014: crom <= 108'o0153_3441_0316_4174_4007_0700_0010_0000_0000;
            12'o2015: crom <= 108'o3217_3441_1603_4174_4007_0700_0000_0000_0000;
            12'o2016: crom <= 108'o2016_3446_1616_4174_4047_0630_2000_0060_0000;
            12'o2017: crom <= 108'o0453_3221_0017_4174_4007_0700_0000_0000_0000;
            12'o2020: crom <= 108'o2020_3444_0303_4174_4047_0630_2000_0060_0000;
            12'o2021: crom <= 108'o3230_3446_1200_4174_4007_0700_0000_0000_0000;
            12'o2022: crom <= 108'o0732_5547_0606_4374_4007_0701_0000_0077_7400;
            12'o2023: crom <= 108'o0732_3547_0606_4374_4007_0701_0000_0077_7400;
            12'o2024: crom <= 108'o2025_0002_0500_4174_4007_0700_0000_0000_0000;
            12'o2025: crom <= 108'o3240_3444_0303_4174_4047_0700_0000_0000_0000;
            12'o2026: crom <= 108'o2027_0002_0500_4174_4007_0700_0000_0000_0000;
            12'o2027: crom <= 108'o0520_3333_0003_4174_4003_4701_1000_0041_0002;
            12'o2030: crom <= 108'o3243_4557_0004_1274_4007_0700_0000_0000_1441;
            12'o2031: crom <= 108'o3241_7441_1717_4174_4007_0700_0000_0000_0000;
            12'o2032: crom <= 108'o2034_5547_0303_4374_4007_0701_0000_0077_7400;
            12'o2033: crom <= 108'o3244_7441_1717_4174_4007_0700_0000_0000_0000;
            12'o2034: crom <= 108'o3042_3442_0400_4174_4007_0700_0010_0000_0000;
            12'o2035: crom <= 108'o2036_2113_0305_4174_4007_0521_4000_0000_0000;
            12'o2036: crom <= 108'o0555_4443_0000_4174_4467_0700_0000_0071_1000;
            12'o2037: crom <= 108'o0724_3221_0004_4174_4007_0700_0000_0000_0000;
            12'o2040: crom <= 108'o0520_3441_1603_4174_4003_4701_0000_0000_0000;
            12'o2041: crom <= 108'o0200_3441_1603_4174_4003_4701_0000_0000_0000;
            12'o2042: crom <= 108'o0520_3444_0303_4174_4043_4701_1000_0041_1777;
            12'o2043: crom <= 108'o1515_3440_0303_1174_4007_0700_0400_0000_1441;
            12'o2044: crom <= 108'o3252_7222_0000_4174_4007_0700_0000_0000_0000;
            12'o2045: crom <= 108'o2046_2222_0000_4174_4007_0511_4000_0000_0000;
            12'o2046: crom <= 108'o0200_7441_0303_4174_4003_4701_0000_0000_0000;
            12'o2047: crom <= 108'o0200_2441_0303_4174_4003_4701_4000_0000_0000;
            12'o2050: crom <= 108'o3254_7333_0003_0174_4007_0700_0400_0000_0000;
            12'o2051: crom <= 108'o3254_2443_0300_0174_4007_0701_4400_0000_0000;
            12'o2052: crom <= 108'o0200_3444_0303_4174_4043_4701_1000_0041_1777;
            12'o2053: crom <= 108'o1515_3440_0303_1174_4007_0700_0400_0000_1441;
            12'o2054: crom <= 108'o0023_3551_1313_4374_0004_1700_0000_0000_2000;
            12'o2055: crom <= 108'o0023_5551_1313_4374_0004_1700_0000_0000_2000;
            12'o2056: crom <= 108'o3400_3333_0005_7174_4001_2700_0400_0000_0241;
            12'o2057: crom <= 108'o0556_3771_0005_4374_0007_0700_0000_0077_7777;
            12'o2060: crom <= 108'o3556_4553_0500_4374_4007_0321_0010_0077_7000;
            12'o2061: crom <= 108'o3556_4553_0400_4374_4007_0321_0010_0077_7000;
            12'o2062: crom <= 108'o3460_4521_0306_4374_4007_0700_0010_0077_7000;
            12'o2063: crom <= 108'o2066_2113_0305_1174_4007_0521_4400_0000_1443;
            12'o2064: crom <= 108'o2062_3771_0003_0276_6007_0700_0000_0000_0000;
            12'o2065: crom <= 108'o2110_3771_0006_0276_6007_0700_0000_0000_0000;
            12'o2066: crom <= 108'o3264_7441_0503_4174_4007_0700_0000_0000_0000;
            12'o2067: crom <= 108'o3264_7441_0303_4174_4007_0700_0000_0000_0000;
            12'o2070: crom <= 108'o2070_4224_0003_4174_4026_7701_1000_0041_1770;
            12'o2071: crom <= 108'o3560_4443_0000_4174_4007_0700_0010_0000_0000;
            12'o2072: crom <= 108'o3267_7221_0003_4174_4007_0700_0000_0000_0000;
            12'o2073: crom <= 108'o3302_3771_0003_7274_4007_0701_0000_0000_0211;
            12'o2074: crom <= 108'o3271_3440_0303_1174_4007_0700_0400_0000_1443;
            12'o2075: crom <= 108'o2074_1111_0503_4174_4007_0700_4000_0000_0000;
            12'o2076: crom <= 108'o2077_0111_0503_4174_4007_0700_0000_0000_0000;
            12'o2077: crom <= 108'o3273_3111_0603_4174_4007_0700_0000_0000_0000;
            12'o2100: crom <= 108'o3277_3333_0003_7174_4007_0700_0400_0000_0211;
            12'o2101: crom <= 108'o2102_1111_0704_4174_4007_0521_4000_0000_0000;
            12'o2102: crom <= 108'o0650_3770_0305_4334_4016_7371_0000_0033_6000;
            12'o2103: crom <= 108'o0546_4223_0000_1174_4007_0700_0400_0000_1443;
            12'o2104: crom <= 108'o3664_0111_0403_4174_4007_0700_0010_0000_0000;
            12'o2105: crom <= 108'o3720_3113_0306_0174_4007_0700_0400_0000_0000;
            12'o2106: crom <= 108'o2107_0111_0703_4174_4007_0700_0000_0000_0000;
            12'o2107: crom <= 108'o2112_0111_0703_4170_4007_0700_0200_0004_0012;
            12'o2110: crom <= 108'o3556_4553_0600_4374_4007_0321_0010_0077_7000;
            12'o2111: crom <= 108'o3556_4553_0600_4374_4007_0321_0010_0004_7777;
            12'o2112: crom <= 108'o3662_4221_0003_4174_4007_0700_0010_0000_0000;
            12'o2113: crom <= 108'o3320_3223_0000_7174_4007_0700_0400_0000_0244;
            12'o2114: crom <= 108'o2106_2113_0604_4174_4007_0521_4000_0000_0000;
            12'o2115: crom <= 108'o3401_3443_0600_4174_4007_0700_0200_0004_0012;
            12'o2116: crom <= 108'o0250_4221_0013_4170_4003_7700_0000_0000_0000;
            12'o2117: crom <= 108'o3311_3771_0003_1276_6007_0701_0000_0000_1441;
            12'o2120: crom <= 108'o3323_3772_0000_7274_4007_0701_0000_0000_0244;
            12'o2121: crom <= 108'o2116_4221_0003_4174_4007_0700_0000_0000_0000;
            12'o2122: crom <= 108'o3451_3771_0003_1276_6007_0701_0010_0000_1444;
            12'o2123: crom <= 108'o0340_3333_0003_4174_4006_5701_1000_0051_0770;
            12'o2124: crom <= 108'o2220_3771_0004_1276_6007_0701_0010_0000_1444;
            12'o2125: crom <= 108'o2220_3333_0004_7174_4007_0700_0410_0000_0250;
            12'o2126: crom <= 108'o2130_3440_0404_1174_4007_0700_0400_0000_1444;
            12'o2127: crom <= 108'o2160_3333_0003_7174_4007_0520_0400_0000_0247;
            12'o2130: crom <= 108'o2154_3333_0006_4174_4007_0520_0010_0000_0000;
            12'o2131: crom <= 108'o0616_4551_0303_4374_0003_7700_0000_0000_0777;
            12'o2132: crom <= 108'o3335_7771_0003_7274_4007_0701_0000_0000_0242;
            12'o2133: crom <= 108'o1050_3771_0005_1276_6007_0622_0000_0000_1443;
            12'o2134: crom <= 108'o1050_4443_0000_4174_4007_0700_0000_0000_0000;
            12'o2135: crom <= 108'o3332_3775_0005_1276_6007_0701_0000_0000_1444;
            12'o2136: crom <= 108'o3665_0551_0505_1274_4007_0700_0010_0000_1444;
            12'o2137: crom <= 108'o0460_0113_0305_1174_4007_0701_0400_0000_1444;
            12'o2140: crom <= 108'o0004_4443_0000_4174_4004_1700_0000_0000_0000;
            12'o2141: crom <= 108'o3334_4551_0404_4374_0007_0700_0000_0037_7777;
            12'o2142: crom <= 108'o3341_3771_0004_1276_6007_0701_0000_0000_1444;
            12'o2143: crom <= 108'o3337_3771_0003_1276_6007_0701_0000_0000_1444;
            12'o2144: crom <= 108'o3340_4551_0303_4374_0007_0700_0000_0037_7777;
            12'o2145: crom <= 108'o3340_3551_0303_4374_0007_0700_0000_0040_0000;
            12'o2146: crom <= 108'o2154_3770_0606_0174_4007_0520_0410_0000_0000;
            12'o2147: crom <= 108'o0260_4221_0013_4170_4007_0700_0000_0000_0000;
            12'o2150: crom <= 108'o2153_7771_0003_1274_4007_0700_0000_0000_1443;
            12'o2151: crom <= 108'o2152_1771_0003_1274_4007_0621_4000_0000_1443;
            12'o2152: crom <= 108'o2153_4571_1204_4374_4007_0700_0000_0040_0000;
            12'o2153: crom <= 108'o3343_3440_0303_1174_4007_0700_0400_0000_1443;
            12'o2154: crom <= 108'o3344_4223_0000_1174_4007_0700_0400_0000_1443;
            12'o2155: crom <= 108'o0001_4443_0000_4174_4004_1700_0000_0000_0000;
            12'o2156: crom <= 108'o3345_4551_0606_4374_4007_0700_0000_0077_7000;
            12'o2157: crom <= 108'o3363_3771_0003_0276_6007_0700_0000_0000_0000;
            12'o2160: crom <= 108'o2170_4221_0006_4170_4007_0700_0000_0000_0000;
            12'o2161: crom <= 108'o2164_3551_0606_4374_0007_0700_0000_0010_0000;
            12'o2162: crom <= 108'o2160_3440_0404_1174_4007_0700_0400_0000_1441;
            12'o2163: crom <= 108'o3347_0111_0704_4174_4007_0700_0000_0000_0000;
            12'o2164: crom <= 108'o3071_4551_0404_4374_0007_0700_0010_0037_7777;
            12'o2165: crom <= 108'o2220_3441_1617_4174_4007_0700_0210_0000_0010;
            12'o2166: crom <= 108'o2162_3770_0303_0174_4007_0520_0400_0000_0000;
            12'o2167: crom <= 108'o2216_1551_0404_6274_4007_0561_4000_0000_0000;
            12'o2170: crom <= 108'o0441_3771_0003_0276_6007_0700_0000_0000_0000;
            12'o2171: crom <= 108'o2174_3551_0606_4374_0007_0700_0000_0020_0000;
            12'o2172: crom <= 108'o2174_3551_0606_4374_0007_0700_0000_0020_0000;
            12'o2173: crom <= 108'o2174_0111_0706_4174_4007_0700_0000_0000_0000;
            12'o2174: crom <= 108'o3460_3771_0003_1276_6007_0701_0010_0000_1443;
            12'o2175: crom <= 108'o3350_4221_0005_4174_4007_0700_0000_0000_0000;
            12'o2176: crom <= 108'o3373_3771_0004_7274_4007_0701_0000_0000_0250;
            12'o2177: crom <= 108'o2200_3333_0006_4174_4007_0520_0000_0000_0000;
            12'o2200: crom <= 108'o2157_3440_0606_1174_4007_0700_0400_0000_1443;
            12'o2201: crom <= 108'o3352_3441_0603_4174_0007_0700_0000_0000_0000;
            12'o2202: crom <= 108'o3374_0111_0704_4174_4007_0700_0000_0000_0000;
            12'o2203: crom <= 108'o3370_3440_0303_0174_4007_0700_0400_0000_0000;
            12'o2204: crom <= 108'o0562_2441_0705_4174_4467_0701_4000_0003_0000;
            12'o2205: crom <= 108'o0260_4221_0013_4170_4467_0700_0000_0005_0000;
            12'o2206: crom <= 108'o3660_4221_0013_4170_4007_0700_0010_0000_0000;
            12'o2207: crom <= 108'o2210_4553_0600_4374_4007_0331_0000_0077_7777;
            12'o2210: crom <= 108'o0637_4221_0003_4174_0007_0700_0000_0000_0000;
            12'o2211: crom <= 108'o2212_4553_0600_4374_4007_0321_0000_0010_0000;
            12'o2212: crom <= 108'o2213_3770_0303_4344_4007_0700_0000_0000_0000;
            12'o2213: crom <= 108'o0637_4221_0003_4174_0007_0700_0000_0000_0000;
            12'o2214: crom <= 108'o2165_0551_0616_4374_4007_0701_0000_0000_0344;
            12'o2215: crom <= 108'o2677_4443_0000_4174_4007_0700_0000_0000_0000;
            12'o2216: crom <= 108'o2217_1111_0703_4174_4007_0700_4000_0000_0000;
            12'o2217: crom <= 108'o3375_0551_0616_4374_4007_0701_0000_0000_0373;
            12'o2220: crom <= 108'o0002_4551_0404_4374_0004_1700_0000_0037_7777;
            12'o2221: crom <= 108'o3377_0551_0303_6274_4007_0700_0000_0000_0000;
            12'o2222: crom <= 108'o0006_4551_0404_4374_0004_1700_0000_0037_7777;
            12'o2223: crom <= 108'o2222_0111_0703_4174_4007_0700_0000_0000_0000;
            12'o2224: crom <= 108'o3660_0115_0505_4174_4007_0700_0010_0000_0000;
            12'o2225: crom <= 108'o0654_3333_0005_4174_4003_1701_0000_0000_0000;
            12'o2226: crom <= 108'o2226_3447_0303_4174_4007_0630_2000_0060_0000;
            12'o2227: crom <= 108'o3403_4551_0303_4374_4007_0700_0000_0000_0777;
            12'o2230: crom <= 108'o2230_3447_0505_4174_4007_0630_2000_0060_0000;
            12'o2231: crom <= 108'o0661_3333_0005_4174_4003_5701_0000_0000_0000;
            12'o2232: crom <= 108'o3423_4443_0000_4174_4007_0700_0000_0000_0000;
            12'o2233: crom <= 108'o0710_3333_0003_4174_4003_5701_0000_0000_0000;
            12'o2234: crom <= 108'o1515_3770_0303_4334_4017_0700_0000_0041_0000;
            12'o2235: crom <= 108'o2234_0111_0703_4174_4007_0700_1000_0051_0700;
            12'o2236: crom <= 108'o3660_3772_0000_1275_5007_0701_0010_0000_1444;
            12'o2237: crom <= 108'o3407_4443_0000_4174_4007_0700_0200_0003_0002;
            12'o2240: crom <= 108'o2275_3771_0003_1276_6007_0701_0010_0000_1441;
            12'o2241: crom <= 108'o0360_3333_0003_4174_4006_5701_0010_0000_0000;
            12'o2242: crom <= 108'o0700_3447_0303_7174_4007_0700_0000_0000_0241;
            12'o2243: crom <= 108'o0006_4443_0000_4174_4004_1700_0000_0000_0000;
            12'o2244: crom <= 108'o0705_4443_0000_4174_4007_0700_0000_0000_0000;
            12'o2245: crom <= 108'o3423_4443_0000_4174_4007_0700_0000_0000_0000;
            12'o2246: crom <= 108'o3417_4751_1203_4374_4007_0700_0010_0000_0002;
            12'o2247: crom <= 108'o0740_3771_0003_4365_5007_0621_0200_0000_0002;
            12'o2250: crom <= 108'o0760_3771_0003_7274_4007_0622_0000_0000_0244;
            12'o2251: crom <= 108'o2252_4251_0303_4374_4007_0700_0000_0000_0077;
            12'o2252: crom <= 108'o3417_0111_0703_7174_4007_0700_0010_0000_0240;
            12'o2253: crom <= 108'o0760_3771_0003_4365_5007_0700_0200_0000_0002;
            12'o2254: crom <= 108'o3421_4551_0303_4374_4007_0700_0000_0000_0077;
            12'o2255: crom <= 108'o3423_4443_0000_4174_4007_0700_0000_0000_0000;
            12'o2256: crom <= 108'o2260_3447_0303_4174_4007_0700_2000_0071_0000;
            12'o2257: crom <= 108'o2256_3551_0303_4370_4007_0700_0000_0000_0200;
            12'o2260: crom <= 108'o2260_3447_0303_4174_4007_0630_2000_0060_0000;
            12'o2261: crom <= 108'o3432_0111_0306_4170_4007_0700_0000_0000_0000;
            12'o2262: crom <= 108'o0002_4443_0000_4174_4004_1700_0000_0000_0000;
            12'o2263: crom <= 108'o0332_4443_0000_7174_4007_0700_0000_0000_0244;
            12'o2264: crom <= 108'o3661_3445_0303_4174_4007_0700_0010_0000_0000;
            12'o2265: crom <= 108'o2266_4553_0300_4374_4007_0331_0000_0000_0001;
            12'o2266: crom <= 108'o0721_3441_0403_4174_4003_1701_0000_0000_0000;
            12'o2267: crom <= 108'o2266_3770_0404_4344_4007_0700_0000_0000_0000;
            12'o2270: crom <= 108'o0754_3333_0004_4174_4003_7530_0000_0000_0000;
            12'o2271: crom <= 108'o0005_4251_0403_4374_4004_1700_0000_0007_7777;
            12'o2272: crom <= 108'o1074_3771_0003_7274_4007_0701_0000_0000_0242;
            12'o2273: crom <= 108'o1074_0551_0703_7274_4007_0701_0000_0000_0242;
            12'o2274: crom <= 108'o0001_3771_0003_1276_6004_1701_0000_0000_1443;
            12'o2275: crom <= 108'o3445_3771_0003_1276_6007_0701_0000_0000_1441;
            12'o2276: crom <= 108'o3076_3333_0003_4174_4217_0701_1010_0073_0500;
            12'o2277: crom <= 108'o0340_3333_0003_4174_4006_5701_1000_0051_0770;
            12'o2300: crom <= 108'o3451_3771_0003_1276_6007_0701_0010_0000_1444;
            12'o2301: crom <= 108'o2241_0113_0404_4174_4007_0701_1000_0077_0000;
            12'o2302: crom <= 108'o3473_3771_0003_1276_6007_0701_0010_0000_1441;
            12'o2303: crom <= 108'o2700_3440_0505_1174_4007_0700_0400_0000_1441;
            12'o2304: crom <= 108'o3453_3441_0503_4174_4217_0700_0000_0000_0600;
            12'o2305: crom <= 108'o3572_0111_0703_4174_4007_0700_0010_0000_0000;
            12'o2306: crom <= 108'o3452_3770_0503_4334_4017_0700_0000_0032_6000;
            12'o2307: crom <= 108'o2356_4221_0003_4174_4007_0700_0000_0000_0000;
            12'o2310: crom <= 108'o3473_3771_0003_1276_6007_0701_0010_0000_1444;
            12'o2311: crom <= 108'o2700_3440_0505_1174_4007_0700_0400_0000_1444;
            12'o2312: crom <= 108'o3466_3440_0303_1174_4007_0700_0400_0000_1443;
            12'o2313: crom <= 108'o2314_3441_0304_4174_4007_0700_0000_0000_0000;
            12'o2314: crom <= 108'o3671_3551_0404_7274_4007_0701_0010_0000_0214;
            12'o2315: crom <= 108'o3465_1111_0503_4174_4007_0700_4000_0000_0000;
            12'o2316: crom <= 108'o3476_0111_1103_4364_4007_0700_0200_0024_1016;
            12'o2317: crom <= 108'o3476_0111_1003_4364_4007_0700_0200_0024_1016;
            12'o2320: crom <= 108'o2716_4443_0000_4174_4467_0700_0000_0001_0000;
            12'o2321: crom <= 108'o2737_4551_0202_4374_0007_0700_0000_0077_7740;
            12'o2322: crom <= 108'o2323_3111_0405_4174_4007_0700_0000_0000_0000;
            12'o2323: crom <= 108'o2324_4553_0300_4374_4007_0331_0000_0004_0000;
            12'o2324: crom <= 108'o2325_5111_0405_4174_4007_0700_0000_0000_0000;
            12'o2325: crom <= 108'o3510_3771_0006_4304_4007_0701_0000_0000_0000;
            12'o2326: crom <= 108'o2327_5111_0406_4174_4007_0700_0000_0000_0000;
            12'o2327: crom <= 108'o2330_4553_0300_4374_4007_0331_0000_0001_0000;
            12'o2330: crom <= 108'o2331_3111_0406_4174_4007_0700_0000_0000_0000;
            12'o2331: crom <= 108'o2332_4553_0300_4374_4007_0331_0000_0003_0000;
            12'o2332: crom <= 108'o3513_3333_0006_4174_4007_0700_0000_0000_0000;
            12'o2333: crom <= 108'o3511_3333_0005_4174_4007_0700_0000_0000_0000;
            12'o2334: crom <= 108'o2336_4551_0303_4374_0007_0321_0000_0010_0000;
            12'o2335: crom <= 108'o3525_4551_1111_4374_0007_0700_0000_0077_0077;
            12'o2336: crom <= 108'o3527_4551_0305_4374_4007_0700_0000_0000_3777;
            12'o2337: crom <= 108'o1400_3111_0311_4174_0477_0700_0000_0000_0000;
            12'o2340: crom <= 108'o2340_3445_0505_4174_4007_0630_2000_0060_0000;
            12'o2341: crom <= 108'o3530_4551_1111_4374_0007_0700_0000_0077_7774;
            12'o2342: crom <= 108'o2342_3445_0303_4174_4007_0630_2000_0060_0000;
            12'o2343: crom <= 108'o3533_3771_0005_7274_4007_0701_0000_0000_0230;
            12'o2344: crom <= 108'o2345_3551_0505_4370_4007_0700_0000_0003_0000;
            12'o2345: crom <= 108'o3535_3333_0005_4174_4257_0700_0000_0000_0000;
            12'o2346: crom <= 108'o2406_3551_1010_4374_0007_0700_0000_0040_0000;
            12'o2347: crom <= 108'o2406_5551_1010_4374_0007_0700_0000_0040_0000;
            12'o2350: crom <= 108'o2350_3447_0505_4174_4007_0630_2000_0060_0000;
            12'o2351: crom <= 108'o3540_4551_0505_4374_4007_0700_0000_0006_3777;
            12'o2352: crom <= 108'o2354_3447_1106_4174_4007_0700_2010_0071_0006;
            12'o2353: crom <= 108'o3614_3443_0300_4174_4007_0700_0200_0003_0012;
            12'o2354: crom <= 108'o2354_3447_0606_4174_4007_0630_2000_0060_0000;
            12'o2355: crom <= 108'o3543_4551_0606_4374_4007_0700_0000_0000_3777;
            12'o2356: crom <= 108'o3564_3333_0003_7174_4007_0700_0400_0000_0301;
            12'o2357: crom <= 108'o2305_3771_0003_7274_4007_0701_0000_0000_0300;
            12'o2360: crom <= 108'o0002_3333_0003_7174_4004_1700_0400_0000_0303;
            12'o2361: crom <= 108'o3566_3771_0003_7274_4007_0701_0000_0000_0302;
            12'o2362: crom <= 108'o2363_3441_0604_4174_4007_0700_0000_0000_0000;
            12'o2363: crom <= 108'o3576_3771_0005_7274_4007_0701_0000_0000_0300;
            12'o2364: crom <= 108'o2365_4221_0014_4174_4007_0700_0000_0000_0000;
            12'o2365: crom <= 108'o2366_4553_0300_4374_4007_0331_0000_0074_0000;
            12'o2366: crom <= 108'o2737_4551_0202_4374_0007_0700_0000_0077_7740;
            12'o2367: crom <= 108'o3605_4551_0305_4374_4007_0700_0000_0000_0177;
            12'o2370: crom <= 108'o2371_5111_0514_4174_0007_0700_0000_0000_0000;
            12'o2371: crom <= 108'o2372_4553_0300_4374_4007_0331_0000_0000_4000;
            12'o2372: crom <= 108'o2373_3111_0514_4174_0007_0700_0000_0000_0000;
            12'o2373: crom <= 108'o2374_4553_0300_4374_4007_0331_0000_0000_0200;
            12'o2374: crom <= 108'o2375_3551_1414_4370_4007_0700_0000_0000_0200;
            12'o2375: crom <= 108'o2376_4553_0300_4374_4007_0331_0000_0000_0400;
            12'o2376: crom <= 108'o2377_5551_1414_4370_4007_0700_0000_0000_0200;
            12'o2377: crom <= 108'o2400_4553_0300_4374_4007_0331_0000_0000_2000;
            12'o2400: crom <= 108'o2401_3111_0514_4170_4007_0700_0000_0000_0000;
            12'o2401: crom <= 108'o0304_4553_0300_4374_4007_0331_0000_0000_1000;
            12'o2402: crom <= 108'o3621_3771_0003_4374_4007_0700_0010_0037_7377;
            12'o2403: crom <= 108'o3616_3771_0005_4374_4247_0700_0000_0000_1001;
            12'o2404: crom <= 108'o2404_1111_0503_4174_4247_0630_6000_0060_1000;
            12'o2405: crom <= 108'o2411_3333_0003_4174_4007_0700_0000_0000_0000;
            12'o2406: crom <= 108'o3621_3771_0003_4374_4007_0700_0010_0037_7377;
            12'o2407: crom <= 108'o3617_3771_0005_4374_4347_0700_0000_0000_1001;
            12'o2410: crom <= 108'o2410_1111_0503_4174_4347_0630_6000_0060_1000;
            12'o2411: crom <= 108'o3620_4223_0000_7174_4007_0700_0400_0000_0424;
            12'o2412: crom <= 108'o3666_4571_1203_4374_4007_0700_0010_0024_1300;
            12'o2413: crom <= 108'o2414_3771_0003_4364_4007_0331_0200_0000_0002;
            12'o2414: crom <= 108'o3642_4221_0004_4174_4007_0700_0000_0000_0000;
            12'o2415: crom <= 108'o3634_3445_0603_4174_4007_0700_0000_0000_0000;
            12'o2416: crom <= 108'o2420_6553_0300_4374_4007_0321_0000_0026_4000;
            12'o2417: crom <= 108'o3641_4521_1205_4074_4007_0700_0000_0000_0000;
            12'o2420: crom <= 108'o0104_4751_1217_4374_4007_0700_0000_0000_0101;
            12'o2421: crom <= 108'o0470_4443_0000_4174_4007_0700_0200_0023_0002;
            12'o2422: crom <= 108'o3642_0111_1504_4174_4007_0700_0000_0000_0000;
            12'o2423: crom <= 108'o2424_4571_1203_4374_4007_0700_0000_0024_1240;
            12'o2424: crom <= 108'o3666_3111_0403_4174_4007_0700_0010_0000_0000;
            12'o2425: crom <= 108'o2426_3771_0016_4364_4007_0700_0200_0000_0002;
            12'o2426: crom <= 108'o3663_0551_1005_4374_4007_0701_0010_0000_0100;
            12'o2427: crom <= 108'o3643_0111_0504_4174_4007_0700_0200_0024_1016;
            12'o2430: crom <= 108'o3644_4557_1606_4374_4007_0701_0000_0000_0774;
            12'o2431: crom <= 108'o0104_4751_1217_4374_4007_0700_0000_0000_0102;
            12'o2432: crom <= 108'o3646_3771_0005_4374_4007_0700_0000_0004_0000;
            12'o2433: crom <= 108'o0004_4443_0000_4174_4004_1700_0000_0000_0000;
            12'o2434: crom <= 108'o0004_5111_0514_4170_4004_1700_0000_0000_0000;
            12'o2435: crom <= 108'o3646_3447_0505_4174_4007_0700_0000_0000_0000;
            12'o2436: crom <= 108'o2456_4443_0000_4174_4137_0700_0010_0000_0000;
            12'o2437: crom <= 108'o0067_4443_0000_4174_4003_7700_0000_0000_0000;
            12'o2440: crom <= 108'o3656_3113_0305_4174_4007_0701_0210_0000_0036;
            12'o2441: crom <= 108'o1027_3771_0005_4364_4003_7700_0200_0000_0002;
            12'o2442: crom <= 108'o2444_3447_0505_4174_4007_0700_2000_0071_0005;
            12'o2443: crom <= 108'o0003_4551_0503_4374_4004_1700_0000_0000_0377;
            12'o2444: crom <= 108'o2444_3447_0505_4174_4007_0630_2000_0060_0000;
            12'o2445: crom <= 108'o0003_4551_0503_4374_4004_1700_0000_0000_0377;
            12'o2446: crom <= 108'o2456_4443_0000_4174_4137_0700_0010_0000_0000;
            12'o2447: crom <= 108'o0227_4443_0000_4174_4003_7700_0000_0000_0000;
            12'o2450: crom <= 108'o3656_3333_0005_4175_5007_0701_0210_0000_0002;
            12'o2451: crom <= 108'o0110_3443_0100_4174_4156_4700_0200_0014_0012;
            12'o2452: crom <= 108'o2454_3445_0505_4174_4007_0700_2000_0071_0005;
            12'o2453: crom <= 108'o3650_4571_1204_4374_4007_0700_0000_0021_1220;
            12'o2454: crom <= 108'o2454_3445_0505_4174_4007_0630_2000_0060_0000;
            12'o2455: crom <= 108'o3650_4571_1204_4374_4007_0700_0000_0021_1220;
            12'o2456: crom <= 108'o3660_1113_0701_4170_4007_0700_4210_0004_0012;
            12'o2457: crom <= 108'o3651_7441_0306_4174_4007_0700_0000_0000_0000;
            12'o2460: crom <= 108'o2462_4553_0200_4374_4007_0321_0000_0000_0020;
            12'o2461: crom <= 108'o2460_4713_1203_7174_4007_0700_0400_0000_0422;
            12'o2462: crom <= 108'o3652_3771_0003_7274_4007_0701_0000_0000_0422;
            12'o2463: crom <= 108'o1055_4443_0000_2174_4006_6700_0000_0000_0000;
            12'o2464: crom <= 108'o2465_0551_0303_2270_4007_0701_0000_0000_0000;
            12'o2465: crom <= 108'o3654_3443_0300_4174_4007_0700_0200_0004_0012;
            12'o2466: crom <= 108'o0001_0551_0403_7274_4124_1701_0000_0000_0422;
            12'o2467: crom <= 108'o3655_0551_0403_7274_4007_0701_0000_0000_0422;
            12'o2470: crom <= 108'o2472_4443_0000_4174_4127_0630_2000_0060_0000;
            12'o2471: crom <= 108'o0001_4443_0000_4174_4004_1700_0000_0000_0000;
            12'o2472: crom <= 108'o2470_4443_0000_4174_4127_0653_0000_0000_0000;
            12'o2473: crom <= 108'o1501_4571_1206_4374_4007_0700_0000_0020_0000;
            12'o2474: crom <= 108'o3670_0111_0704_4170_4007_0700_0210_0023_1016;
            12'o2475: crom <= 108'o0005_4443_0000_4174_4107_0700_0000_0000_0074;
            12'o2476: crom <= 108'o0117_3443_0100_4174_4007_0700_0200_0014_0012;
            12'o2477: crom <= 108'o2500_4571_1203_4374_4007_0700_0000_0024_1200;
            12'o2500: crom <= 108'o3666_3551_0303_4370_4007_0700_0010_0020_0000;
            12'o2501: crom <= 108'o2716_3771_0002_4365_5617_0700_0200_0000_0002;
            12'o2502: crom <= 108'o3700_3333_0012_4174_4437_0700_0000_0000_0000;
            12'o2503: crom <= 108'o0002_3771_0004_7274_4004_1701_0000_0000_0212;
            12'o2504: crom <= 108'o2746_3333_0000_4175_5007_0701_0210_0000_0002;
            12'o2505: crom <= 108'o2746_3333_0002_4175_5007_0701_0210_0000_0002;
            12'o2506: crom <= 108'o3701_3333_0001_4175_5007_0701_0200_0000_0002;
            12'o2507: crom <= 108'o2510_3333_0003_4175_5007_0701_0200_0000_0002;
            12'o2510: crom <= 108'o2746_3333_0003_7174_4007_0700_0410_0000_0211;
            12'o2511: crom <= 108'o2746_3333_0003_4175_5007_0701_0210_0000_0002;
            12'o2512: crom <= 108'o2511_3771_0003_7274_4007_0701_0000_0000_0212;
            12'o2513: crom <= 108'o3702_3333_0005_4175_5007_0701_0200_0000_0002;
            12'o2514: crom <= 108'o2746_3333_0006_4175_5007_0701_0210_0000_0002;
            12'o2515: crom <= 108'o2746_3333_0010_4175_5007_0701_0210_0000_0002;
            12'o2516: crom <= 108'o3703_3333_0007_4175_5007_0701_0200_0000_0002;
            12'o2517: crom <= 108'o3704_3333_0011_4175_5007_0701_0200_0000_0002;
            12'o2520: crom <= 108'o2746_3333_0012_4175_5007_0701_0210_0000_0002;
            12'o2521: crom <= 108'o2746_3333_0014_4175_5007_0701_0210_0000_0002;
            12'o2522: crom <= 108'o3705_3333_0013_4175_5007_0701_0200_0000_0002;
            12'o2523: crom <= 108'o3706_3333_0015_4175_5007_0701_0200_0000_0002;
            12'o2524: crom <= 108'o2746_3333_0016_4175_5007_0701_0210_0000_0002;
            12'o2525: crom <= 108'o2746_3771_0003_7274_4007_0701_0010_0000_0210;
            12'o2526: crom <= 108'o2525_3333_0017_4175_5007_0701_0200_0000_0002;
            12'o2527: crom <= 108'o3707_3333_0003_4175_5007_0701_0200_0000_0002;
            12'o2530: crom <= 108'o3727_3771_0013_4370_4007_0700_0000_0040_0002;
            12'o2531: crom <= 108'o0100_3440_0303_0174_4156_4700_0400_0000_0000;
            12'o2532: crom <= 108'o2533_3551_0606_4374_0007_0700_0000_0001_0000;
            12'o2533: crom <= 108'o3732_4551_0606_4374_0007_0700_0000_0041_1000;
            12'o2534: crom <= 108'o2534_3447_0505_4174_4007_0630_2000_0060_0000;
            12'o2535: crom <= 108'o3734_4251_0505_4374_4007_0700_0000_0000_0777;
            12'o2536: crom <= 108'o2540_3333_0006_4174_4007_0520_0000_0000_0000;
            12'o2537: crom <= 108'o3774_3447_0504_4174_4007_0700_0000_0000_0000;
            12'o2540: crom <= 108'o2544_3771_0004_7274_4007_0622_0000_0000_0423;
            12'o2541: crom <= 108'o2542_3771_0004_7274_4007_0622_0000_0000_0424;
            12'o2542: crom <= 108'o1130_0113_0405_4174_4007_0700_0200_0024_1016;
            12'o2543: crom <= 108'o3735_0551_1103_4374_4007_0701_0000_0000_0540;
            12'o2544: crom <= 108'o1130_0113_0405_4174_4007_0700_0200_0024_1016;
            12'o2545: crom <= 108'o3735_0551_1003_4374_4007_0701_0000_0000_0540;
            12'o2546: crom <= 108'o2672_4553_1300_4374_4007_0321_0000_0001_0000;
            12'o2547: crom <= 108'o0602_3445_0303_4174_4007_0630_2000_0060_0000;
            12'o2550: crom <= 108'o3772_4443_0000_4174_4007_0700_0010_0000_0000;
            12'o2551: crom <= 108'o0030_4443_0000_2174_4006_6700_0000_0000_0000;
            12'o2552: crom <= 108'o2672_4553_1300_4374_4007_0321_0000_0001_0000;
            12'o2553: crom <= 108'o2555_4251_0304_4374_4007_0700_0000_0000_3777;
            12'o2554: crom <= 108'o2552_4553_0300_4374_4007_0321_0000_0000_0077;
            12'o2555: crom <= 108'o2622_3441_0403_4174_4007_0700_0010_0000_0000;
            12'o2556: crom <= 108'o2551_3771_0002_4365_5217_0700_0200_0000_0002;
            12'o2557: crom <= 108'o2560_3551_0303_7274_4007_0701_0000_0000_0220;
            12'o2560: crom <= 108'o3075_4443_0000_4174_4007_0700_0210_0001_0002;
            12'o2561: crom <= 108'o3772_4443_0000_4174_4007_0700_0010_0000_0000;
            12'o2562: crom <= 108'o2562_3445_0404_4174_4007_0630_2000_0060_0000;
            12'o2563: crom <= 108'o1040_3333_0006_4174_4007_0520_0000_0000_0000;
            12'o2564: crom <= 108'o2562_4443_0000_4174_4007_0700_2000_0071_0007;
            12'o2565: crom <= 108'o1134_4553_0300_4374_4007_0321_0000_0000_0077;
            12'o2566: crom <= 108'o2600_3333_0003_7174_4007_0700_0400_0000_0426;
            12'o2567: crom <= 108'o2570_4251_0505_4374_4007_0370_0000_0000_0777;
            12'o2570: crom <= 108'o1000_4551_0303_4374_0007_0700_0000_0027_7000;
            12'o2571: crom <= 108'o2672_4553_1300_4374_4007_0321_0000_0001_0000;
            12'o2572: crom <= 108'o3745_3551_0606_4374_4007_0700_0000_0002_0000;
            12'o2573: crom <= 108'o2574_4553_0600_4374_4007_0321_0000_0003_0000;
            12'o2574: crom <= 108'o2672_4553_1300_4374_4007_0321_0000_0001_0000;
            12'o2575: crom <= 108'o2603_3551_0303_7274_4007_0701_0000_0000_0220;
            12'o2576: crom <= 108'o2604_3551_0303_4370_4007_0700_0000_0000_0001;
            12'o2577: crom <= 108'o2604_4553_0300_4374_4007_0331_0000_0000_0001;
            12'o2600: crom <= 108'o3561_3771_0003_7274_4117_0701_0010_0000_0301;
            12'o2601: crom <= 108'o0104_4751_1217_4374_4007_0700_0000_0000_0001;
            12'o2602: crom <= 108'o1133_3771_0003_7274_4007_0701_0000_0000_0426;
            12'o2603: crom <= 108'o3075_4443_0000_4174_4007_0700_0210_0001_0002;
            12'o2604: crom <= 108'o2575_3551_0606_4374_0007_0700_0000_0004_0000;
            12'o2605: crom <= 108'o2575_5551_1313_4374_0007_0700_0000_0002_0000;
            12'o2606: crom <= 108'o2623_3771_0005_4365_5007_0700_0200_0000_0002;
            12'o2607: crom <= 108'o2610_4553_1300_4374_4007_0331_0000_0040_0000;
            12'o2610: crom <= 108'o2612_3441_0403_4174_4007_0700_2000_0071_0007;
            12'o2611: crom <= 108'o3753_3771_0003_7274_4007_0701_0000_0000_0210;
            12'o2612: crom <= 108'o2612_3445_0303_4174_4007_0630_2000_0060_0000;
            12'o2613: crom <= 108'o3746_4551_0303_4374_0007_0700_0000_0000_0003;
            12'o2614: crom <= 108'o2615_3551_0606_4374_0007_0700_0000_0000_2000;
            12'o2615: crom <= 108'o3752_4551_0606_4370_4007_0700_0000_0000_0777;
            12'o2616: crom <= 108'o2617_3551_0606_4374_4007_0700_0000_0004_0000;
            12'o2617: crom <= 108'o2620_4553_1300_4374_4147_0321_0000_0000_4000;
            12'o2620: crom <= 108'o3762_3551_0606_4374_4007_0700_0000_0002_0000;
            12'o2621: crom <= 108'o3762_3333_0006_4174_4007_0700_0000_0000_0000;
            12'o2622: crom <= 108'o3772_0551_0303_7274_4007_0701_0010_0000_0216;
            12'o2623: crom <= 108'o2627_0111_0703_4174_4007_0700_0200_0004_0012;
            12'o2624: crom <= 108'o0002_4551_0303_7274_4004_1701_0000_0000_0217;
            12'o2625: crom <= 108'o2672_4553_1300_4374_4007_0321_0000_0001_0000;
            12'o2626: crom <= 108'o2624_4553_0300_4374_4007_0321_0000_0077_0000;
            12'o2627: crom <= 108'o2701_3771_0001_4361_5007_0700_0200_0000_0002;
            12'o2630: crom <= 108'o2632_4553_0300_4374_4007_0321_0000_0030_0000;
            12'o2631: crom <= 108'o2672_4553_1300_4374_4007_0321_0000_0001_0000;
            12'o2632: crom <= 108'o2634_4553_0300_4374_4007_0321_0000_0010_0000;
            12'o2633: crom <= 108'o2672_4553_1300_4374_4007_0321_0000_0001_0000;
            12'o2634: crom <= 108'o2636_4553_0300_4374_4007_0321_0000_0020_0000;
            12'o2635: crom <= 108'o0002_4443_0000_4174_4004_1700_0000_0000_0000;
            12'o2636: crom <= 108'o0003_4443_0000_4174_4004_1700_0000_0000_0000;
            12'o2637: crom <= 108'o0001_4443_0000_4174_4004_1700_0000_0000_0000;
            12'o2640: crom <= 108'o0004_3771_0003_4365_5004_1700_0200_0000_0002;
            12'o2641: crom <= 108'o2672_4553_1300_4374_4007_0321_0000_0001_0000;
            12'o2642: crom <= 108'o0007_4443_0000_4174_4004_1700_0000_0000_0000;
            12'o2643: crom <= 108'o3773_7441_1303_4174_4007_0700_0000_0000_0000;
            12'o2644: crom <= 108'o0007_4443_0000_4174_4004_1700_0000_0000_0000;
            12'o2645: crom <= 108'o0002_4443_0000_4174_4004_1700_0000_0000_0000;
            12'o2646: crom <= 108'o2650_1553_0500_4374_4007_0532_4000_0000_0340;
            12'o2647: crom <= 108'o3775_0111_1104_4174_4007_0700_0200_0024_1016;
            12'o2650: crom <= 108'o2652_1553_0500_4374_4007_0532_4000_0000_0400;
            12'o2651: crom <= 108'o2652_0551_0404_4374_4007_0701_0000_0000_0600;
            12'o2652: crom <= 108'o3775_0111_1004_4174_4007_0700_0200_0024_1016;
            12'o2653: crom <= 108'o2647_0551_0404_4374_4007_0701_0000_0000_0220;
            12'o2654: crom <= 108'o2656_3333_0004_4174_4007_0530_0000_0000_0000;
            12'o2655: crom <= 108'o2654_3770_0404_4344_4007_0700_0000_0000_0000;
            12'o2656: crom <= 108'o2672_4553_1300_4374_4007_0321_0000_0001_0000;
            12'o2657: crom <= 108'o1435_5551_1313_4374_4007_0700_0000_0002_4000;
            12'o2660: crom <= 108'o2661_3551_1313_4374_0007_0700_0000_0000_4000;
            12'o2661: crom <= 108'o2662_4553_0400_4374_4007_0331_0000_0004_0000;
            12'o2662: crom <= 108'o2663_3551_0606_4374_0007_0700_0000_0002_0000;
            12'o2663: crom <= 108'o2664_4553_0400_4374_4007_0331_0000_0010_0000;
            12'o2664: crom <= 108'o1500_3551_1313_4374_0007_0700_0000_0002_0000;
            12'o2665: crom <= 108'o2666_4553_0600_4374_4007_0321_0000_0001_0000;
            12'o2666: crom <= 108'o2656_3551_0606_4374_0007_0700_0000_0010_0000;
            12'o2667: crom <= 108'o2607_4443_0000_4174_4007_0700_0000_0000_0000;
            12'o2670: crom <= 108'o1510_3771_0005_4354_4007_0700_0010_0000_0000;
            12'o2671: crom <= 108'o1502_4551_0505_4374_0007_0700_0000_0040_1237;
            12'o2672: crom <= 108'o0104_4751_1217_4374_4007_0700_0000_0000_0100;
            12'o2673: crom <= 108'o2674_3771_0003_7274_4007_0611_0000_0000_0210;
            12'o2674: crom <= 108'o2676_4553_0300_4374_4007_0321_0000_0010_0000;
            12'o2675: crom <= 108'o1511_3771_0003_7274_4007_0701_0000_0000_0425;
            12'o2676: crom <= 108'o1100_4443_0000_4174_4007_0700_0000_0000_0000;
            12'o2677: crom <= 108'o2700_1111_0701_4170_4007_0700_4000_0000_0000;
            12'o2700: crom <= 108'o1100_3333_0013_4174_4003_5701_0000_0000_0000;
            12'o2701: crom <= 108'o2714_3333_0005_4174_4467_0700_0000_0001_0004;
            12'o2702: crom <= 108'o1512_0551_1103_4374_4007_0701_0000_0000_0500;
            12'o2703: crom <= 108'o0770_3551_1313_4374_0007_0700_0000_0001_0000;
            12'o2704: crom <= 108'o1564_3333_0006_4175_5007_0701_0210_0000_0002;
            12'o2705: crom <= 108'o2706_4553_1000_4374_4007_0321_0000_0040_0000;
            12'o2706: crom <= 108'o2712_4521_1205_4074_4007_0700_0000_0000_0000;
            12'o2707: crom <= 108'o1513_3741_0105_4074_4007_0700_0000_0000_0000;
            12'o2710: crom <= 108'o1500_3441_0603_4174_4003_7700_0200_0003_0001;
            12'o2711: crom <= 108'o2703_1111_0701_4174_4007_0700_4000_0000_0000;
            12'o2712: crom <= 108'o1564_3333_0005_4175_5007_0701_0210_0000_0002;
            12'o2713: crom <= 108'o1563_3333_0001_4175_5007_0701_0200_0000_0002;
            12'o2714: crom <= 108'o0305_5551_1313_4374_4007_0700_0000_0001_0000;
            12'o2715: crom <= 108'o0435_4521_1203_4074_4007_0700_0000_0000_0000;
            12'o2716: crom <= 108'o0371_4713_1202_7174_4007_0700_0400_0000_0422;
            12'o2717: crom <= 108'o1044_0551_1504_0274_4407_0311_0200_0003_0712;
            12'o2720: crom <= 108'o0220_4443_0000_4174_4463_7700_0000_0001_2000;
            12'o2721: crom <= 108'o2722_3771_0005_4365_5007_0700_0200_0000_0002;
            12'o2722: crom <= 108'o1144_0551_0404_4374_4407_0311_0000_0077_7777;
            12'o2723: crom <= 108'o0220_3333_0005_4175_5003_7701_0200_0000_0002;
            12'o2724: crom <= 108'o2720_3333_0005_4175_5007_0701_0200_0000_0002;
            12'o2725: crom <= 108'o1146_0551_0404_4374_4407_0311_0000_0077_7777;
            12'o2726: crom <= 108'o1150_3771_0005_0276_6007_0521_0000_0000_0000;
            12'o2727: crom <= 108'o0764_3440_0505_0174_4467_0700_0400_0005_0000;
            12'o2730: crom <= 108'o2731_3443_0300_4174_4007_0700_0200_0003_0012;
            12'o2731: crom <= 108'o2732_3333_0005_4175_5007_0701_0200_0000_0002;
            12'o2732: crom <= 108'o1400_0551_0301_4370_4007_0701_0000_0000_0001;
            12'o2733: crom <= 108'o0130_3770_0304_4344_4007_0700_0000_0000_0000;
            12'o2734: crom <= 108'o2735_3770_0505_4344_4007_0700_0000_0000_0000;
            12'o2735: crom <= 108'o2736_3443_0500_4174_4007_0700_0200_0004_0012;
            12'o2736: crom <= 108'o0274_3771_0005_4365_5007_0700_0200_0000_0002;
            12'o2737: crom <= 108'o1156_4751_1204_4374_4007_0700_0000_0000_0424;
            12'o2740: crom <= 108'o2741_0111_1105_4174_4007_0700_0000_0000_0000;
            12'o2741: crom <= 108'o2742_4521_1203_4074_4007_0700_0000_0000_0000;
            12'o2742: crom <= 108'o1164_4553_0300_4374_4007_0321_0000_0000_0600;
            12'o2743: crom <= 108'o2744_3771_0003_4365_5007_0700_0200_0000_0002;
            12'o2744: crom <= 108'o0764_3333_0003_4174_4467_0700_0000_0000_0404;
            12'o2745: crom <= 108'o0001_5551_0303_4374_0004_1700_0000_0000_0600;
            12'o2746: crom <= 108'o0002_0111_0704_4170_4004_1700_0200_0023_1016;
            12'o2747: crom <= 108'o2750_4551_0202_4374_0007_0700_0000_0077_7740;
            12'o2750: crom <= 108'o2751_3333_0002_4175_5007_0701_0200_0000_0002;
            12'o2751: crom <= 108'o2501_0111_0703_4170_4007_0700_0200_0004_0012;
            12'o2752: crom <= 108'o1170_3111_0503_4170_4007_0700_0000_0000_0000;
            12'o2753: crom <= 108'o1174_3770_0303_4174_0007_0520_0000_0000_0000;
            12'o2754: crom <= 108'o0021_3772_0000_0275_5007_0700_2000_0071_0043;
            12'o2755: crom <= 108'o1200_5113_0412_4174_4007_0621_0000_0000_0000;
            12'o2756: crom <= 108'o2757_3441_0316_4174_4007_0700_0000_0000_0000;
            12'o2757: crom <= 108'o0031_3771_0006_0276_6007_0700_2000_0071_0043;
            12'o2760: crom <= 108'o1204_3770_0303_4174_0007_0520_0000_0000_0000;
            12'o2761: crom <= 108'o2762_4117_0004_4174_4007_0700_0000_0000_0000;
            12'o2762: crom <= 108'o0120_3441_0405_4174_4007_0350_0000_0000_0000;
            12'o2763: crom <= 108'o0410_3227_0004_1174_4007_0700_0400_0000_1442;
            12'o2764: crom <= 108'o0410_3777_0016_1276_6007_0701_0000_0000_1441;
            12'o2765: crom <= 108'o0543_0111_1604_4174_4007_0700_0000_0000_0000;
            12'o2766: crom <= 108'o1210_3770_0404_0174_4007_0520_0400_0000_0000;
            12'o2767: crom <= 108'o2770_3772_0000_1275_5007_0701_0000_0000_1442;
            12'o2770: crom <= 108'o2771_7003_0000_1174_4007_0700_0400_0000_1442;
            12'o2771: crom <= 108'o2772_3772_0000_1275_5007_0701_0000_0000_1443;
            12'o2772: crom <= 108'o2773_7003_0000_1174_4007_0700_0400_0000_1443;
            12'o2773: crom <= 108'o1212_3741_0103_4074_4007_0520_0000_0000_0000;
            12'o2774: crom <= 108'o2775_4221_0004_4174_4007_0700_0000_0000_0000;
            12'o2775: crom <= 108'o2776_3442_0500_4174_4007_0700_2000_0071_0043;
            12'o2776: crom <= 108'o0563_3447_0606_4174_4007_0700_0000_0000_0000;
            12'o2777: crom <= 108'o2677_4443_0000_4174_4467_0700_0000_0003_0000;
            12'o3000: crom <= 108'o3001_3446_0606_4174_4007_0700_0000_0000_0000;
            12'o3001: crom <= 108'o0122_4226_0004_4174_4007_0630_2000_0060_0000;
            12'o3002: crom <= 108'o0122_3446_1200_4174_4007_0630_2000_0060_0000;
            12'o3003: crom <= 108'o1214_3772_0000_0275_5007_0520_0000_0000_0000;
            12'o3004: crom <= 108'o3005_3771_0003_0276_6007_0700_0000_0000_0000;
            12'o3005: crom <= 108'o3006_3772_0000_1275_5007_0701_0000_0000_1441;
            12'o3006: crom <= 108'o0160_3333_0003_4174_4007_0621_0000_0000_0000;
            12'o3007: crom <= 108'o3010_3221_0004_4174_4007_0700_0000_0000_0000;
            12'o3010: crom <= 108'o0330_3333_0003_4174_4007_0520_0000_0000_0000;
            12'o3011: crom <= 108'o1224_3447_0305_4174_4007_0421_0000_0000_0000;
            12'o3012: crom <= 108'o3013_3662_0000_4374_0007_0700_0000_0060_0000;
            12'o3013: crom <= 108'o3014_2222_0000_4174_4007_0700_4000_0000_0000;
            12'o3014: crom <= 108'o3016_2446_0505_4174_4047_0700_0040_0000_0000;
            12'o3015: crom <= 108'o3016_4751_1217_4374_4007_0700_0000_0000_0004;
            12'o3016: crom <= 108'o3017_3221_0006_0174_4007_0700_0000_0000_0000;
            12'o3017: crom <= 108'o0054_3777_0003_0274_4007_0520_0000_0000_0000;
            12'o3020: crom <= 108'o0354_4552_0000_1275_5007_0701_0000_0000_1442;
            12'o3021: crom <= 108'o3022_0002_1600_4174_4007_0700_0000_0000_0000;
            12'o3022: crom <= 108'o1242_4003_0000_1174_4007_0700_0400_0000_1440;
            12'o3023: crom <= 108'o0551_4552_0000_1275_5007_0701_0000_0000_1443;
            12'o3024: crom <= 108'o0056_3333_0017_4174_4003_5701_0000_0000_0000;
            12'o3025: crom <= 108'o3026_1772_0000_0274_4007_0701_0040_0000_0000;
            12'o3026: crom <= 108'o1244_3223_0000_0174_4007_0621_0400_0000_0000;
            12'o3027: crom <= 108'o3032_4113_1600_1174_4007_0700_0400_0000_1441;
            12'o3030: crom <= 108'o3031_3551_1616_4374_0007_0700_0000_0040_0000;
            12'o3031: crom <= 108'o3032_3440_1616_1174_4007_0700_0400_0000_1441;
            12'o3032: crom <= 108'o1246_3333_0003_4174_4007_0520_0000_0000_0000;
            12'o3033: crom <= 108'o3034_0111_0503_4174_4007_0700_0040_0000_0000;
            12'o3034: crom <= 108'o3035_0002_0600_4174_4007_0700_0000_0000_0000;
            12'o3035: crom <= 108'o3036_0111_0503_4174_4007_0700_0040_0000_0000;
            12'o3036: crom <= 108'o0355_3333_0017_4174_4003_5701_0000_0000_0000;
            12'o3037: crom <= 108'o3040_2444_0303_4174_4047_0700_0040_0000_0000;
            12'o3040: crom <= 108'o1250_0113_0303_1174_4007_0521_0400_0000_1442;
            12'o3041: crom <= 108'o0100_7003_0000_1174_4156_4700_0400_0000_1443;
            12'o3042: crom <= 108'o0001_3446_0303_4174_4044_1700_0000_0000_0000;
            12'o3043: crom <= 108'o1252_3333_0003_4174_4007_0520_0000_0000_0000;
            12'o3044: crom <= 108'o3045_3771_0004_4374_4007_0700_0000_0010_0000;
            12'o3045: crom <= 108'o1256_3333_0005_4174_4007_0520_0000_0000_0000;
            12'o3046: crom <= 108'o1256_3551_0404_4374_4007_0700_0000_0004_0000;
            12'o3047: crom <= 108'o3050_3447_0303_4174_4007_0700_0000_0000_0000;
            12'o3050: crom <= 108'o3051_3447_0505_4174_4007_0700_0000_0000_0000;
            12'o3051: crom <= 108'o3052_3447_0505_4174_4007_0700_0000_0000_0000;
            12'o3052: crom <= 108'o1260_1114_0503_4174_4067_0630_6000_0060_0000;
            12'o3053: crom <= 108'o1262_3447_0303_4174_4007_0520_0000_0000_0000;
            12'o3054: crom <= 108'o3055_3444_0303_4174_4007_0700_0000_0000_0000;
            12'o3055: crom <= 108'o3056_4002_1200_4174_4007_0700_0000_0000_0000;
            12'o3056: crom <= 108'o0014_3333_0004_4174_4000_1701_0000_0000_0000;
            12'o3057: crom <= 108'o1266_0115_0503_4174_4007_0630_2040_0060_0000;
            12'o3060: crom <= 108'o3061_1772_0000_1274_4007_0701_4000_0000_1443;
            12'o3061: crom <= 108'o1270_4003_0000_1174_4007_0621_0400_0000_1443;
            12'o3062: crom <= 108'o1272_4003_0000_1174_4007_0621_0400_0000_1442;
            12'o3063: crom <= 108'o1274_4003_0000_1174_4007_0621_0400_0000_1441;
            12'o3064: crom <= 108'o1272_4003_0000_1174_4007_0700_0400_0000_1442;
            12'o3065: crom <= 108'o1274_4003_0000_1174_4007_0700_0400_0000_1441;
            12'o3066: crom <= 108'o0024_3440_0303_0174_4004_1700_0400_0000_0000;
            12'o3067: crom <= 108'o3070_4551_0404_4374_0007_0700_0000_0037_7777;
            12'o3070: crom <= 108'o1276_2441_0404_4174_4007_0621_4000_0000_0000;
            12'o3071: crom <= 108'o1300_2441_0404_4174_4007_0621_4000_0000_0000;
            12'o3072: crom <= 108'o3073_3443_0400_4174_4007_0701_1000_0077_0000;
            12'o3073: crom <= 108'o0264_3771_0004_0276_6007_0700_0000_0000_0000;
            12'o3074: crom <= 108'o3075_0111_0703_4170_4007_0700_0200_0003_0002;
            12'o3075: crom <= 108'o0004_3333_0003_4175_5004_1701_0200_0000_0002;
            12'o3076: crom <= 108'o0070_4443_0000_2174_4006_6700_0000_0000_0000;
            12'o3077: crom <= 108'o0070_4443_0000_2174_4466_6700_0000_0003_0000;
            12'o3100: crom <= 108'o3076_3771_0003_4361_5217_0700_0200_0000_0502;
            12'o3101: crom <= 108'o0001_4551_1205_4365_5004_1700_0200_0000_0002;
            12'o3102: crom <= 108'o0002_4257_0503_4374_4004_1701_0000_0000_0376;
            12'o3103: crom <= 108'o3104_4221_0005_4174_0007_0700_1000_0031_0220;
            12'o3104: crom <= 108'o3105_3447_0505_4174_4007_0700_1020_0041_0010;
            12'o3105: crom <= 108'o3106_3333_0003_4174_4007_0700_1000_0031_7770;
            12'o3106: crom <= 108'o3107_4222_0000_4174_4007_0700_0000_0000_0000;
            12'o3107: crom <= 108'o3110_4224_0003_4174_4027_0700_1020_0041_0010;
            12'o3110: crom <= 108'o3111_4224_0003_4174_4027_0700_0000_0000_0000;
            12'o3111: crom <= 108'o0002_4001_0503_4174_4004_1700_0000_0000_0000;
            12'o3112: crom <= 108'o3113_3447_1200_4174_4007_0700_0200_0003_0002;
            12'o3113: crom <= 108'o0002_3333_0003_4175_5004_1701_0200_0000_0002;
            12'o3114: crom <= 108'o3115_4222_0000_4174_4007_0700_0000_0000_0000;
            12'o3115: crom <= 108'o3116_4224_0000_4174_4027_0700_1020_0041_0010;
            12'o3116: crom <= 108'o3117_4224_0000_4174_4027_0700_0000_0000_0000;
            12'o3117: crom <= 108'o3120_3333_0003_4174_4007_0701_1000_0073_0000;
            12'o3120: crom <= 108'o3121_4443_0000_4174_4007_0700_1000_0051_0770;
            12'o3121: crom <= 108'o3122_4002_1200_4174_4007_0700_1000_0031_0000;
            12'o3122: crom <= 108'o3123_3444_0404_4174_4007_0700_1020_0041_0010;
            12'o3123: crom <= 108'o3124_7221_0003_4174_4007_0700_0000_0000_0000;
            12'o3124: crom <= 108'o3125_4111_0503_4174_4007_0700_0000_0000_0000;
            12'o3125: crom <= 108'o3126_4001_0404_4174_4007_0700_0000_0000_0000;
            12'o3126: crom <= 108'o3112_3111_0403_4174_4007_0700_0000_0000_0000;
            12'o3127: crom <= 108'o1302_3770_0304_4344_4007_0700_2000_0071_0011;
            12'o3130: crom <= 108'o3131_3771_0004_4374_0007_0700_0000_0000_0000;
            12'o3131: crom <= 108'o3132_3333_0004_7174_4007_0700_0400_0000_0221;
            12'o3132: crom <= 108'o3133_4557_0305_4374_4007_0701_0000_0000_7700;
            12'o3133: crom <= 108'o3134_3770_0505_4344_4007_0700_2000_0071_0003;
            12'o3134: crom <= 108'o1304_4221_0005_4174_0007_0700_0000_0000_0000;
            12'o3135: crom <= 108'o3136_3772_0000_4370_4007_0700_0000_0000_0044;
            12'o3136: crom <= 108'o3137_1662_0000_7274_4007_0701_4000_0000_0221;
            12'o3137: crom <= 108'o3140_3771_0005_7274_4007_0701_0000_0000_0222;
            12'o3140: crom <= 108'o0664_4443_0000_4174_4007_0700_2000_0071_0042;
            12'o3141: crom <= 108'o3142_3771_0003_4374_4007_0700_0000_0077_7777;
            12'o3142: crom <= 108'o1310_0661_0005_7274_4007_0622_0000_0000_0224;
            12'o3143: crom <= 108'o1312_3333_0003_4174_4007_0421_0000_0000_0000;
            12'o3144: crom <= 108'o1312_0551_0303_7274_4007_0701_0000_0000_0226;
            12'o3145: crom <= 108'o3146_3441_0306_4174_4007_0700_2000_0071_0043;
            12'o3146: crom <= 108'o0062_3772_0000_7274_4007_0701_0000_0000_0222;
            12'o3147: crom <= 108'o3150_2555_0303_4374_4007_0701_4000_0000_0044;
            12'o3150: crom <= 108'o3151_3770_0303_4344_4007_0700_2000_0071_0011;
            12'o3151: crom <= 108'o1314_3771_0003_4370_4007_0700_0000_0000_0000;
            12'o3152: crom <= 108'o1400_3113_0305_0174_4007_0700_0400_0000_0000;
            12'o3153: crom <= 108'o1316_3770_0604_4344_4007_0700_0000_0000_0000;
            12'o3154: crom <= 108'o3155_2112_0306_4174_4007_0700_4000_0000_0000;
            12'o3155: crom <= 108'o3156_0001_0705_4174_4007_0700_0000_0000_0000;
            12'o3156: crom <= 108'o3157_3770_0505_4344_0007_0700_0000_0000_0000;
            12'o3157: crom <= 108'o3160_0551_0505_0274_4407_0701_0000_0000_0000;
            12'o3160: crom <= 108'o0002_3771_0013_4370_4004_1700_0000_0000_0001;
            12'o3161: crom <= 108'o1320_2113_0506_4174_4007_0331_4000_0000_0000;
            12'o3162: crom <= 108'o1322_3223_0000_4174_4007_0671_0200_0000_0002;
            12'o3163: crom <= 108'o1320_3772_0000_4365_5007_0700_0200_0000_0002;
            12'o3164: crom <= 108'o3165_3223_0000_4174_4007_0701_0200_0000_0002;
            12'o3165: crom <= 108'o1330_2113_0603_4174_4007_0521_4000_0000_0000;
            12'o3166: crom <= 108'o3163_0111_0704_4170_4007_0700_0200_0004_0712;
            12'o3167: crom <= 108'o3170_3770_0303_4344_4007_0700_0000_0000_0000;
            12'o3170: crom <= 108'o3171_3771_0003_7270_4007_0701_0000_0000_0214;
            12'o3171: crom <= 108'o1100_3440_0303_0174_4007_0700_0400_0000_0000;
            12'o3172: crom <= 108'o3173_3441_0503_4174_4007_0700_2000_0041_2000;
            12'o3173: crom <= 108'o3174_3441_0405_4174_4007_0700_2000_0020_0000;
            12'o3174: crom <= 108'o1332_3333_0003_4174_4007_0520_1000_0041_2000;
            12'o3175: crom <= 108'o1336_4222_0000_4174_4007_0630_2000_0060_0000;
            12'o3176: crom <= 108'o0163_3442_0300_4174_4007_0700_2000_0071_0033;
            12'o3177: crom <= 108'o3200_3441_0403_4174_4007_0700_1000_0041_0002;
            12'o3200: crom <= 108'o0420_3446_0303_4174_4003_4701_1000_0041_1600;
            12'o3201: crom <= 108'o3203_3441_0304_4174_4007_0700_1000_0031_0200;
            12'o3202: crom <= 108'o3203_2441_0304_4174_4007_0700_5000_0031_0200;
            12'o3203: crom <= 108'o1346_3445_0506_4174_4007_0520_0000_0000_0000;
            12'o3204: crom <= 108'o1363_4222_0000_4174_4007_0700_0000_0000_0000;
            12'o3205: crom <= 108'o1362_3446_0303_4174_4047_0700_2000_0071_0006;
            12'o3206: crom <= 108'o3207_4222_0000_0174_4007_0700_0000_0000_0000;
            12'o3207: crom <= 108'o1364_3771_0003_0276_6007_0520_1000_0040_2000;
            12'o3210: crom <= 108'o1366_4443_0000_4174_4007_0630_2000_0060_0000;
            12'o3211: crom <= 108'o1514_4221_0013_4174_4003_7700_0200_0003_0001;
            12'o3212: crom <= 108'o1637_2441_0303_4174_4007_0700_0040_0000_0000;
            12'o3213: crom <= 108'o2006_3777_0005_0274_4007_0521_2000_0020_2000;
            12'o3214: crom <= 108'o3220_0002_0400_4174_4007_0700_0000_0000_0000;
            12'o3215: crom <= 108'o3216_3442_0400_4174_4007_0700_2000_0020_0000;
            12'o3216: crom <= 108'o2014_3333_0016_4174_4007_0700_1000_0041_2000;
            12'o3217: crom <= 108'o3220_0002_0600_4174_4007_0700_0000_0000_0000;
            12'o3220: crom <= 108'o3221_0116_0503_4174_4047_0700_0040_0000_0000;
            12'o3221: crom <= 108'o0433_3444_0303_4174_4046_2700_0000_0000_0000;
            12'o3222: crom <= 108'o3223_3444_0303_4174_4047_0700_1000_0041_1777;
            12'o3223: crom <= 108'o3224_3444_0303_4174_4047_0700_1000_0041_1777;
            12'o3224: crom <= 108'o2027_3002_1700_4170_4007_0700_0000_0000_0000;
            12'o3225: crom <= 108'o3226_3444_1616_4174_4067_0700_0000_0000_0000;
            12'o3226: crom <= 108'o0472_3446_1616_4174_4047_0630_2000_0060_0000;
            12'o3227: crom <= 108'o0001_3446_1616_4174_4044_1700_0000_0000_0000;
            12'o3230: crom <= 108'o3231_4662_0000_4374_0007_0700_0000_0007_7777;
            12'o3231: crom <= 108'o3232_3221_0005_4174_4007_0700_0000_0000_0000;
            12'o3232: crom <= 108'o0623_4557_0006_1274_4007_0700_0000_0000_1441;
            12'o3233: crom <= 108'o3234_3227_0004_4174_4007_0700_2000_0011_0000;
            12'o3234: crom <= 108'o2022_3777_0006_0274_4007_0521_1000_0040_2000;
            12'o3235: crom <= 108'o1012_0111_1604_4174_4007_0700_0000_0000_0000;
            12'o3236: crom <= 108'o3237_3447_0705_4174_4007_0700_0000_0000_0000;
            12'o3237: crom <= 108'o2024_4553_1700_4374_4007_0321_0000_0020_0000;
            12'o3240: crom <= 108'o2026_4553_1700_4374_4007_0321_0000_0010_0000;
            12'o3241: crom <= 108'o3242_2441_0606_4174_4007_0700_4000_0000_0000;
            12'o3242: crom <= 108'o2030_2331_0005_1174_4007_0521_0040_0000_1441;
            12'o3243: crom <= 108'o2032_3777_0003_0274_4007_0521_1000_0030_2000;
            12'o3244: crom <= 108'o3245_3547_0303_4374_4007_0701_0000_0077_7400;
            12'o3245: crom <= 108'o3246_2442_0400_4174_4007_0700_4000_0000_0000;
            12'o3246: crom <= 108'o2035_2446_0303_4174_4047_0700_0040_0000_0000;
            12'o3247: crom <= 108'o0513_3444_1616_4174_4046_2700_0000_0000_0000;
            12'o3250: crom <= 108'o1515_4113_0400_1174_4007_0700_0400_0000_1441;
            12'o3251: crom <= 108'o2042_3223_0000_4174_4007_0621_0000_0000_0000;
            12'o3252: crom <= 108'o2046_4221_0013_4174_4007_0700_0000_0000_0000;
            12'o3253: crom <= 108'o2050_4221_0013_4174_4007_0700_0000_0000_0000;
            12'o3254: crom <= 108'o0100_4113_0400_1174_4156_4700_0400_0000_1441;
            12'o3255: crom <= 108'o2052_3223_0000_4174_4007_0621_0000_0000_0000;
            12'o3256: crom <= 108'o0002_4553_1300_4374_4004_1321_0000_0000_2000;
            12'o3257: crom <= 108'o3260_3111_0605_4174_0417_0700_0000_0000_0000;
            12'o3260: crom <= 108'o3261_3333_0005_4174_4217_0700_0000_0000_0500;
            12'o3261: crom <= 108'o3262_3333_0003_7174_4007_0700_0400_0000_0240;
            12'o3262: crom <= 108'o0170_4443_0000_2174_4006_6700_0000_0000_0000;
            12'o3263: crom <= 108'o3262_3771_0005_4361_5217_0700_0200_0000_0502;
            12'o3264: crom <= 108'o0574_3333_0003_7174_4003_7700_0400_0000_0242;
            12'o3265: crom <= 108'o3266_3333_0005_4174_4007_0700_1000_0041_6020;
            12'o3266: crom <= 108'o2070_4222_0000_4174_4006_7701_1000_0041_1770;
            12'o3267: crom <= 108'o0507_4113_0312_7174_4007_0700_0400_0000_0243;
            12'o3270: crom <= 108'o2074_3771_0005_1276_6007_0522_0000_0000_1443;
            12'o3271: crom <= 108'o3272_7771_0003_7274_4007_0701_0000_0000_0242;
            12'o3272: crom <= 108'o2076_3333_0005_4174_4007_0520_0000_0000_0000;
            12'o3273: crom <= 108'o1515_4221_0013_4170_4007_0700_0000_0000_0000;
            12'o3274: crom <= 108'o2100_3440_0303_1174_4007_0670_0400_0000_1441;
            12'o3275: crom <= 108'o2104_3440_0303_1174_4007_0700_0400_0000_1443;
            12'o3276: crom <= 108'o3274_0111_0703_4170_4007_0700_0000_0000_0000;
            12'o3277: crom <= 108'o3300_3333_0005_7174_4007_0700_0400_0000_0213;
            12'o3300: crom <= 108'o3301_3333_0004_7174_4007_0700_0400_0000_0212;
            12'o3301: crom <= 108'o2071_3333_0006_7174_4007_0700_0400_0000_0214;
            12'o3302: crom <= 108'o3303_3771_0005_7274_4007_0701_0000_0000_0213;
            12'o3303: crom <= 108'o3304_3771_0004_7274_4007_0701_0000_0000_0212;
            12'o3304: crom <= 108'o3274_3771_0006_7274_4007_0701_0000_0000_0214;
            12'o3305: crom <= 108'o3306_0111_0704_4174_4007_0700_0000_0000_0000;
            12'o3306: crom <= 108'o0540_3771_0013_4370_4007_0700_0000_0000_0003;
            12'o3307: crom <= 108'o3310_3113_0406_0174_4007_0700_0400_0000_0000;
            12'o3310: crom <= 108'o0252_4221_0013_4170_4007_0700_0000_0000_0000;
            12'o3311: crom <= 108'o1020_3333_0006_4174_4007_0520_0000_0000_0000;
            12'o3312: crom <= 108'o3313_3440_0606_0174_4007_0700_0400_0000_0000;
            12'o3313: crom <= 108'o3314_3771_0013_4370_4007_0700_0000_0000_0010;
            12'o3314: crom <= 108'o1030_3333_0004_4174_4007_0520_0000_0000_0000;
            12'o3315: crom <= 108'o3316_4111_1203_7174_4007_0700_0000_0000_0245;
            12'o3316: crom <= 108'o3317_4551_1205_7274_4007_0700_0000_0000_0245;
            12'o3317: crom <= 108'o3320_2111_0503_4174_4007_0700_4000_0000_0000;
            12'o3320: crom <= 108'o3321_1111_0704_4174_4007_0700_4000_0000_0000;
            12'o3321: crom <= 108'o3322_1111_0706_4174_4007_0700_4000_0000_0000;
            12'o3322: crom <= 108'o2116_3333_0003_4174_4007_0621_0000_0000_0000;
            12'o3323: crom <= 108'o3324_3771_0013_4370_4007_0700_0000_0000_0012;
            12'o3324: crom <= 108'o1030_3223_0000_7174_4007_0700_0400_0000_0245;
            12'o3325: crom <= 108'o3326_3333_0003_7174_4007_0700_0400_0000_0243;
            12'o3326: crom <= 108'o3327_3771_0003_0276_6007_0700_0000_0000_0000;
            12'o3327: crom <= 108'o2124_4521_0306_4374_4007_0700_0000_0077_7000;
            12'o3330: crom <= 108'o0460_7333_0003_7174_4007_0700_0400_0000_0242;
            12'o3331: crom <= 108'o2134_4553_0500_4374_4007_0321_0000_0076_0000;
            12'o3332: crom <= 108'o2136_3445_0505_1174_4007_0700_0000_0000_1444;
            12'o3333: crom <= 108'o0002_3440_0505_1174_4004_1700_0400_0000_1443;
            12'o3334: crom <= 108'o0004_0111_0705_4174_4004_1700_0000_0000_0000;
            12'o3335: crom <= 108'o3336_3111_0306_4174_4007_0700_0000_0000_0000;
            12'o3336: crom <= 108'o2143_1111_0701_4170_4007_0700_4000_0000_0000;
            12'o3337: crom <= 108'o2144_3771_0005_1276_6007_0522_0000_0000_1443;
            12'o3340: crom <= 108'o2146_3440_0303_1174_4007_0700_0400_0000_1444;
            12'o3341: crom <= 108'o3342_4551_0404_4374_0007_0700_0000_0037_7777;
            12'o3342: crom <= 108'o2150_2441_0404_1174_4007_0621_4000_0000_1443;
            12'o3343: crom <= 108'o2143_3440_0404_1174_4007_0700_0400_0000_1444;
            12'o3344: crom <= 108'o0001_4223_0000_1174_4004_1700_0400_0000_1444;
            12'o3345: crom <= 108'o3346_3771_0004_1276_6007_0701_0000_0000_1441;
            12'o3346: crom <= 108'o2125_3771_0003_0276_6007_0700_2000_0071_0024;
            12'o3347: crom <= 108'o2164_3551_0606_4374_0007_0700_0000_0004_0000;
            12'o3350: crom <= 108'o3351_3441_0605_4170_4007_0700_0000_0000_0000;
            12'o3351: crom <= 108'o2176_1111_0305_4174_4007_0421_4000_0000_0000;
            12'o3352: crom <= 108'o3353_3440_0303_1174_4007_0700_0400_0000_1443;
            12'o3353: crom <= 108'o3354_3771_0003_7274_4007_0701_0000_0000_0240;
            12'o3354: crom <= 108'o3355_0111_0703_4174_4007_0700_0200_0004_0012;
            12'o3355: crom <= 108'o3356_3771_0016_4365_5007_0700_0200_0000_0002;
            12'o3356: crom <= 108'o3357_3771_0013_4370_4007_0700_0000_0000_0012;
            12'o3357: crom <= 108'o3360_2113_0507_7174_4007_0701_4400_0000_0242;
            12'o3360: crom <= 108'o3361_3441_1603_7174_4007_0700_0000_0000_0242;
            12'o3361: crom <= 108'o0640_0551_0705_7274_4007_0521_0000_0000_0242;
            12'o3362: crom <= 108'o3360_3440_0505_1174_4007_0700_0400_0000_1443;
            12'o3363: crom <= 108'o3372_3771_0004_1276_6007_0701_0000_0000_1441;
            12'o3364: crom <= 108'o0636_0551_0503_7274_4003_7701_0000_0000_0241;
            12'o3365: crom <= 108'o3366_3771_0003_7274_4007_0701_0000_0000_0247;
            12'o3366: crom <= 108'o3367_3771_0004_7274_4007_0701_0000_0000_0250;
            12'o3367: crom <= 108'o2202_4553_0500_4374_4007_0321_0000_0004_0000;
            12'o3370: crom <= 108'o3371_3440_0404_1174_4007_0700_0400_0000_1441;
            12'o3371: crom <= 108'o3372_3440_0505_1174_4007_0700_0400_0000_1443;
            12'o3372: crom <= 108'o2204_1111_0706_4174_4007_0531_4000_0000_0000;
            12'o3373: crom <= 108'o1505_3771_0003_7274_4007_0701_0000_0000_0247;
            12'o3374: crom <= 108'o2203_5551_0505_4374_0007_0700_0000_0004_0000;
            12'o3375: crom <= 108'o3376_3333_0016_4174_4007_0700_0200_0000_0010;
            12'o3376: crom <= 108'o2220_1551_0303_6274_4007_0522_4000_0000_0000;
            12'o3377: crom <= 108'o3400_3333_0017_4174_4007_0700_0200_0000_0010;
            12'o3400: crom <= 108'o2222_0551_0404_6274_4007_0561_0000_0000_0000;
            12'o3401: crom <= 108'o3402_4221_0013_4170_4007_0700_0000_0000_0000;
            12'o3402: crom <= 108'o2224_3770_0605_4344_4007_0700_0000_0000_0000;
            12'o3403: crom <= 108'o2230_3447_0305_4174_4007_0700_2000_0071_0002;
            12'o3404: crom <= 108'o3405_7441_0605_4174_4007_0700_1000_0071_0010;
            12'o3405: crom <= 108'o3406_3441_0603_4174_4007_0701_1000_0043_0000;
            12'o3406: crom <= 108'o2234_4553_0500_4374_4007_0321_0000_0003_0000;
            12'o3407: crom <= 108'o3410_3223_0000_4174_4007_0701_0200_0000_0002;
            12'o3410: crom <= 108'o3423_3440_0303_1174_4007_0700_0400_0000_1444;
            12'o3411: crom <= 108'o0705_4251_0303_4374_4007_0700_0000_0007_7777;
            12'o3412: crom <= 108'o3413_3771_0005_1276_6007_0701_0000_0000_1443;
            12'o3413: crom <= 108'o3414_3443_0500_4174_4007_0700_0200_0003_0012;
            12'o3414: crom <= 108'o3415_3771_0005_1276_6007_0701_0000_0000_1444;
            12'o3415: crom <= 108'o2246_3333_0005_4175_5007_0701_0200_0000_0002;
            12'o3416: crom <= 108'o0007_3440_0606_0174_4004_1700_0400_0000_0000;
            12'o3417: crom <= 108'o3420_0551_0303_7274_4007_0701_0000_0000_0240;
            12'o3420: crom <= 108'o0001_3443_0300_4174_4004_1700_0200_0004_0012;
            12'o3421: crom <= 108'o3422_0115_0703_4174_4007_0700_0000_0000_0000;
            12'o3422: crom <= 108'o3424_3333_0003_4174_4007_0701_2000_0007_0000;
            12'o3423: crom <= 108'o3424_4443_0000_4174_4007_0700_2000_0071_0000;
            12'o3424: crom <= 108'o3425_3333_0006_4174_4007_0701_1000_0073_0000;
            12'o3425: crom <= 108'o3426_4443_0000_4174_4007_0700_1000_0051_0030;
            12'o3426: crom <= 108'o3427_4443_0000_4174_4007_0700_1000_0040_0000;
            12'o3427: crom <= 108'o3430_4443_0000_4174_4007_0700_1000_0041_0010;
            12'o3430: crom <= 108'o3431_3777_0003_4334_4057_0700_2000_0041_0000;
            12'o3431: crom <= 108'o2256_4251_0303_4374_4007_0630_0000_0000_0170;
            12'o3432: crom <= 108'o3433_3770_0303_4334_4017_0700_0000_0041_0000;
            12'o3433: crom <= 108'o3434_4551_0606_4374_0007_0700_0000_0070_0000;
            12'o3434: crom <= 108'o3435_4551_0303_4374_4007_0700_0000_0003_0000;
            12'o3435: crom <= 108'o3436_3111_0306_4174_0007_0700_0000_0000_0000;
            12'o3436: crom <= 108'o2115_3440_0606_0174_4007_0700_0400_0000_0000;
            12'o3437: crom <= 108'o2262_0113_0703_1174_4007_0521_0400_0000_1443;
            12'o3440: crom <= 108'o3441_0551_0303_7274_4007_0700_0000_0000_0241;
            12'o3441: crom <= 108'o0004_4553_0300_7274_4004_1622_0000_0000_0243;
            12'o3442: crom <= 108'o3443_0551_0303_7274_4007_0701_0000_0000_0241;
            12'o3443: crom <= 108'o2264_3333_0003_4174_4007_0700_0200_0004_0012;
            12'o3444: crom <= 108'o2272_3770_0303_1174_4007_0520_0400_0000_1443;
            12'o3445: crom <= 108'o0231_3770_0305_4334_4016_7701_0000_0033_6000;
            12'o3446: crom <= 108'o3447_0111_0703_4170_4007_0700_0000_0000_0000;
            12'o3447: crom <= 108'o2276_3440_0303_1174_4007_0700_0400_0000_1441;
            12'o3450: crom <= 108'o2300_3441_0304_4174_4007_0700_0000_0000_0000;
            12'o3451: crom <= 108'o2304_3770_0305_4334_4016_7701_0000_0033_6000;
            12'o3452: crom <= 108'o3453_0111_0703_4170_4217_0700_0000_0000_0600;
            12'o3453: crom <= 108'o0230_3440_0303_1174_4006_6701_1400_0073_1444;
            12'o3454: crom <= 108'o3455_3771_0003_4361_5217_0700_0200_0000_0602;
            12'o3455: crom <= 108'o0230_4443_0000_2174_4006_6700_0000_0000_0000;
            12'o3456: crom <= 108'o3457_3771_0003_4365_5007_0700_0200_0000_0002;
            12'o3457: crom <= 108'o0010_3333_0003_7174_4004_1700_0400_0000_0244;
            12'o3460: crom <= 108'o0001_4551_0303_4374_0004_1700_0000_0000_0777;
            12'o3461: crom <= 108'o3462_3771_0003_7274_4007_0701_0000_0000_0214;
            12'o3462: crom <= 108'o2310_0113_0703_0174_4007_0701_0400_0000_0000;
            12'o3463: crom <= 108'o3464_1771_0003_7274_4007_0701_4000_0000_0242;
            12'o3464: crom <= 108'o2312_3771_0005_1276_6007_0522_0000_0000_1443;
            12'o3465: crom <= 108'o2700_3440_0303_1174_4007_0700_0400_0000_1443;
            12'o3466: crom <= 108'o3470_0111_0503_4174_4007_0700_0000_0000_0000;
            12'o3467: crom <= 108'o3470_1771_0003_7274_4007_0701_4000_0000_0242;
            12'o3470: crom <= 108'o3471_3551_0303_7274_4007_0701_0000_0000_0214;
            12'o3471: crom <= 108'o2700_3440_0303_0174_4007_0700_0400_0000_0000;
            12'o3472: crom <= 108'o3464_7771_0003_7274_4007_0701_0000_0000_0242;
            12'o3473: crom <= 108'o0001_3770_0305_4334_4014_1700_0000_0043_6000;
            12'o3474: crom <= 108'o3475_3741_0104_4074_4007_0700_0000_0000_0000;
            12'o3475: crom <= 108'o2316_3333_0004_7174_4007_0340_0400_0000_0425;
            12'o3476: crom <= 108'o3477_3771_0002_4365_5617_0700_0200_0000_0002;
            12'o3477: crom <= 108'o2320_4553_0200_4374_4007_0321_0000_0070_0000;
            12'o3500: crom <= 108'o3501_4251_0505_4374_4007_0700_0000_0000_7770;
            12'o3501: crom <= 108'o0260_4113_0305_4174_4007_0330_0000_0000_0000;
            12'o3502: crom <= 108'o0136_4251_0505_4374_4007_0700_0000_0000_7770;
            12'o3503: crom <= 108'o3504_5551_0505_4370_4007_0700_0000_0000_0007;
            12'o3504: crom <= 108'o3505_4551_0304_4374_4007_0700_0000_0000_0007;
            12'o3505: crom <= 108'o3506_3111_0405_4174_4007_0700_0000_0000_0000;
            12'o3506: crom <= 108'o3507_4551_0304_4374_4007_0700_0000_0000_7760;
            12'o3507: crom <= 108'o2322_4553_0300_4374_4007_0331_0000_0010_0000;
            12'o3510: crom <= 108'o2326_4553_0300_4374_4007_0331_0000_0002_0000;
            12'o3511: crom <= 108'o3512_3333_0005_4174_4257_0700_0000_0000_0000;
            12'o3512: crom <= 108'o1400_3333_0005_7174_4007_0700_0400_0000_0230;
            12'o3513: crom <= 108'o3514_3333_0006_4174_4237_0700_0000_0000_0000;
            12'o3514: crom <= 108'o3515_5551_0606_4370_4007_0700_0000_0000_2000;
            12'o3515: crom <= 108'o2333_3333_0006_4174_4237_0700_0000_0000_0000;
            12'o3516: crom <= 108'o3517_3770_0505_4344_0007_0700_0000_0000_0000;
            12'o3517: crom <= 108'o3520_4551_0505_4374_0007_0700_0000_0000_7760;
            12'o3520: crom <= 108'o3521_4551_0505_4370_4007_0700_0000_0000_0007;
            12'o3521: crom <= 108'o3522_3771_0004_4304_4007_0701_0000_0000_0000;
            12'o3522: crom <= 108'o3523_4251_0404_4374_4007_0700_0000_0000_7770;
            12'o3523: crom <= 108'o3613_3111_0405_4174_4007_0700_0000_0000_0000;
            12'o3524: crom <= 108'o2334_3771_0003_4365_5007_0521_0200_0000_0002;
            12'o3525: crom <= 108'o3526_4551_0303_4374_0007_0700_0000_0050_7700;
            12'o3526: crom <= 108'o2336_4553_0300_4374_4007_0321_0000_0010_0000;
            12'o3527: crom <= 108'o2340_4221_0005_4174_0007_0700_2000_0071_0007;
            12'o3530: crom <= 108'o3531_4221_0011_4170_4007_0700_0000_0000_0000;
            12'o3531: crom <= 108'o3532_3111_0511_4174_4007_0700_0000_0000_0000;
            12'o3532: crom <= 108'o2406_3111_0311_4174_0477_0700_0000_0000_0000;
            12'o3533: crom <= 108'o3534_4551_0505_4370_4007_0700_0000_0074_7777;
            12'o3534: crom <= 108'o2344_4553_0300_4374_4007_0321_0000_0000_0020;
            12'o3535: crom <= 108'o3536_3333_0005_7174_4007_0700_0400_0000_0230;
            12'o3536: crom <= 108'o3537_3441_0310_4174_4007_0700_0000_0000_0000;
            12'o3537: crom <= 108'o2346_4553_1000_4374_4007_0321_0000_0000_0040;
            12'o3540: crom <= 108'o3613_4221_0005_4174_0007_0700_0000_0000_0000;
            12'o3541: crom <= 108'o3542_4551_1105_4374_0007_0700_0000_0050_7700;
            12'o3542: crom <= 108'o2354_3447_1106_4174_4007_0700_2000_0071_0006;
            12'o3543: crom <= 108'o0001_3441_0605_4170_4004_1700_0000_0000_0000;
            12'o3544: crom <= 108'o3545_3771_0003_4365_5007_0700_0200_0000_0002;
            12'o3545: crom <= 108'o1400_3333_0003_7174_4007_0700_0400_0000_0215;
            12'o3546: crom <= 108'o3547_3771_0003_4365_5007_0700_0200_0000_0002;
            12'o3547: crom <= 108'o1400_3333_0003_7174_4007_0700_0400_0000_0216;
            12'o3550: crom <= 108'o3551_3771_0003_4365_5007_0700_0200_0000_0002;
            12'o3551: crom <= 108'o1400_3333_0003_7174_4007_0700_0400_0000_0220;
            12'o3552: crom <= 108'o3553_3771_0003_4365_5007_0700_0200_0000_0002;
            12'o3553: crom <= 108'o1400_3333_0003_7174_4007_0700_0400_0000_0217;
            12'o3554: crom <= 108'o3555_3771_0003_4365_5007_0700_0200_0000_0002;
            12'o3555: crom <= 108'o1400_3333_0003_7174_4007_0700_0400_0000_0227;
            12'o3556: crom <= 108'o2737_4551_0202_4374_0007_0700_0000_0077_7740;
            12'o3557: crom <= 108'o0004_4443_0000_4174_4004_1700_0000_0000_0000;
            12'o3560: crom <= 108'o3561_3771_0003_7274_4117_0701_0000_0000_0301;
            12'o3561: crom <= 108'o3562_4751_1205_4374_4007_0700_0000_0001_0000;
            12'o3562: crom <= 108'o3563_0111_0503_4174_4007_0700_0000_0000_0000;
            12'o3563: crom <= 108'o2356_3770_0303_4174_0007_0520_0000_0000_0000;
            12'o3564: crom <= 108'o3565_3771_0003_7274_4007_0701_0000_0000_0303;
            12'o3565: crom <= 108'o2360_1111_0503_4174_4007_0421_4000_0000_0000;
            12'o3566: crom <= 108'o3567_3771_0005_4304_4007_0701_0000_0000_0000;
            12'o3567: crom <= 108'o3570_3551_0505_4374_4007_0700_0000_0000_0040;
            12'o3570: crom <= 108'o2360_3333_0005_4174_4237_0700_0000_0000_0000;
            12'o3571: crom <= 108'o1114_3771_0003_4365_5007_0700_0200_0000_0002;
            12'o3572: crom <= 108'o0002_3333_0003_7174_4004_1700_0400_0000_0300;
            12'o3573: crom <= 108'o3574_4451_1204_4324_4007_0700_0000_0000_0000;
            12'o3574: crom <= 108'o3575_4451_1206_4324_4007_0700_0000_0000_0000;
            12'o3575: crom <= 108'o2362_6113_0405_4174_4007_0621_0000_0000_0000;
            12'o3576: crom <= 108'o1120_0551_0404_7274_4007_0671_0000_0000_0301;
            12'o3577: crom <= 108'o3600_3333_0005_4175_5007_0701_0200_0000_0002;
            12'o3600: crom <= 108'o3601_0111_0702_4170_4007_0700_0200_0003_0012;
            12'o3601: crom <= 108'o1400_3333_0004_4175_5007_0701_0200_0000_0002;
            12'o3602: crom <= 108'o3603_3771_0003_4365_5007_0700_0200_0000_0002;
            12'o3603: crom <= 108'o3604_3333_0003_7174_4007_0700_0400_0000_0302;
            12'o3604: crom <= 108'o1400_3333_0003_7174_4007_0700_0400_0000_0303;
            12'o3605: crom <= 108'o3606_3770_0505_4344_0007_0700_0000_0000_0000;
            12'o3606: crom <= 108'o2370_4553_0300_4374_4007_0331_0000_0002_0000;
            12'o3607: crom <= 108'o3610_3770_1416_4344_4007_0700_0000_0000_0000;
            12'o3610: crom <= 108'o3611_2441_0716_4170_4007_0700_4000_0000_0000;
            12'o3611: crom <= 108'o3612_4111_1416_4174_4007_0700_0000_0000_0000;
            12'o3612: crom <= 108'o0010_7443_1600_4174_4434_1700_0000_0000_0000;
            12'o3613: crom <= 108'o3614_3443_0300_4174_4007_0700_0200_0003_0012;
            12'o3614: crom <= 108'o1400_3333_0005_4175_5007_0701_0200_0000_0002;
            12'o3615: crom <= 108'o2402_4221_0003_4174_4007_0700_0000_0000_0000;
            12'o3616: crom <= 108'o2404_3333_0003_4174_4247_0700_0000_0000_1000;
            12'o3617: crom <= 108'o2410_3333_0003_4174_4347_0700_0000_0000_1000;
            12'o3620: crom <= 108'o1400_4223_0000_7174_4007_0700_0400_0000_0423;
            12'o3621: crom <= 108'o0001_4443_0000_4174_4004_1700_2000_0071_0375;
            12'o3622: crom <= 108'o3631_4751_1206_4374_4007_0700_0000_0000_0001;
            12'o3623: crom <= 108'o3631_4751_1206_4374_4007_0700_0000_0000_0002;
            12'o3624: crom <= 108'o3631_4751_1206_4374_4007_0700_0000_0000_0003;
            12'o3625: crom <= 108'o3631_4751_1206_4374_4007_0700_0000_0000_0004;
            12'o3626: crom <= 108'o3631_4751_1206_4374_4007_0700_0000_0000_0005;
            12'o3627: crom <= 108'o3631_4751_1206_4374_4007_0700_0000_0000_0006;
            12'o3630: crom <= 108'o3631_4751_1206_4374_4007_0700_0000_0000_0007;
            12'o3631: crom <= 108'o3632_4251_1403_4374_4007_0700_0000_0007_7577;
            12'o3632: crom <= 108'o3633_7443_0300_4174_4437_0700_0000_0000_0000;
            12'o3633: crom <= 108'o2412_4223_0000_4364_4277_0700_0200_0000_0010;
            12'o3634: crom <= 108'o3635_0551_0303_4370_4007_0701_0000_0000_0040;
            12'o3635: crom <= 108'o3636_0111_1003_4174_4007_0700_0000_0000_0000;
            12'o3636: crom <= 108'o3637_3443_0300_4174_4007_0700_0200_0024_1016;
            12'o3637: crom <= 108'o3640_3771_0003_4365_5007_0701_0200_0020_0012;
            12'o3640: crom <= 108'o2416_6553_0300_4374_4007_0321_0000_0025_4340;
            12'o3641: crom <= 108'o0060_4223_0000_4174_4467_0700_0000_0000_0004;
            12'o3642: crom <= 108'o2422_3445_0303_4174_4007_0530_0000_0000_0000;
            12'o3643: crom <= 108'o2430_3771_0005_4365_5007_0331_0200_0000_0002;
            12'o3644: crom <= 108'o3645_3447_0606_4174_4007_0700_0000_0000_0000;
            12'o3645: crom <= 108'o3637_0111_0605_4174_4007_0700_0200_0024_0012;
            12'o3646: crom <= 108'o2434_4113_0514_4174_4007_0330_0000_0000_0000;
            12'o3647: crom <= 108'o2446_3441_0603_4174_4007_0700_0000_0000_0000;
            12'o3650: crom <= 108'o2450_3113_0304_4174_4007_0701_0200_0000_0036;
            12'o3651: crom <= 108'o2460_4553_0600_4374_4007_0321_0000_0070_0000;
            12'o3652: crom <= 108'o3653_3333_0002_4174_4217_0700_0000_0000_0000;
            12'o3653: crom <= 108'o2464_4553_0200_4374_4007_0321_0000_0000_0017;
            12'o3654: crom <= 108'o0001_3771_0003_4365_5124_1700_0200_0000_0002;
            12'o3655: crom <= 108'o0001_4221_0003_4174_0124_1700_0000_0000_0000;
            12'o3656: crom <= 108'o1124_3771_0016_4354_4007_0650_2000_0071_0200;
            12'o3657: crom <= 108'o2470_4443_0000_4174_4007_0650_2000_0071_0777;
            12'o3660: crom <= 108'o0001_3771_0003_4365_5004_1700_0200_0000_0002;
            12'o3661: crom <= 108'o0001_3771_0004_4365_5004_1700_0200_0000_0002;
            12'o3662: crom <= 108'o0001_3772_0000_4365_5004_1700_0200_0000_0002;
            12'o3663: crom <= 108'o0001_4221_0004_4174_0004_1700_0000_0000_0000;
            12'o3664: crom <= 108'o0001_0111_0703_4174_4004_1700_0000_0000_0000;
            12'o3665: crom <= 108'o0001_3445_0505_4174_4004_1700_0000_0000_0000;
            12'o3666: crom <= 108'o0001_3443_0300_4174_4004_1701_0200_0000_0036;
            12'o3667: crom <= 108'o0004_3333_0005_4175_5004_1701_0200_0000_0002;
            12'o3670: crom <= 108'o0001_3333_0001_4175_5004_1701_0200_0000_0002;
            12'o3671: crom <= 108'o0001_3440_0404_0174_4004_1700_0400_0000_0000;
            12'o3672: crom <= 108'o1515_3771_0003_4365_5007_0700_0200_0000_0002;
            12'o3673: crom <= 108'o1516_3771_0003_0276_6007_0700_0000_0000_0000;
            12'o3674: crom <= 108'o2474_3333_0017_4175_5007_0701_0200_0000_0002;
            12'o3675: crom <= 108'o2502_3771_0004_7274_4007_0422_0000_0000_0227;
            12'o3676: crom <= 108'o3677_3771_0004_4354_4007_0700_0000_0000_0000;
            12'o3677: crom <= 108'o0010_3333_0004_7174_4004_1700_0400_0000_0210;
            12'o3700: crom <= 108'o2504_3333_0004_4174_4007_0700_0200_0021_1016;
            12'o3701: crom <= 108'o2505_0111_0704_4170_4007_0700_0200_0023_1016;
            12'o3702: crom <= 108'o2514_0111_0704_4170_4007_0700_0200_0023_1016;
            12'o3703: crom <= 108'o2515_0111_0704_4170_4007_0700_0200_0023_1016;
            12'o3704: crom <= 108'o2520_0111_0704_4170_4007_0700_0200_0023_1016;
            12'o3705: crom <= 108'o2521_0111_0704_4170_4007_0700_0200_0023_1016;
            12'o3706: crom <= 108'o2524_0111_0704_4170_4007_0700_0200_0023_1016;
            12'o3707: crom <= 108'o3710_3771_0003_7274_4007_0701_0000_0000_0211;
            12'o3710: crom <= 108'o3711_3771_0004_7274_4007_0701_0000_0000_0210;
            12'o3711: crom <= 108'o3712_3443_0400_4174_4007_0700_0200_0000_0010;
            12'o3712: crom <= 108'o0006_3771_0004_7274_4004_1701_0000_0000_0212;
            12'o3713: crom <= 108'o3714_3771_0006_4354_4007_0700_0000_0000_0000;
            12'o3714: crom <= 108'o3715_4551_0606_4374_0007_0700_0000_0040_0000;
            12'o3715: crom <= 108'o3716_3333_0006_7174_4007_0700_0400_0000_0210;
            12'o3716: crom <= 108'o3717_3771_0005_7274_4007_0701_0000_0000_0230;
            12'o3717: crom <= 108'o2530_4553_0500_4374_4007_0331_0000_0003_0000;
            12'o3720: crom <= 108'o3721_3333_0006_7174_4007_0700_0400_0000_0214;
            12'o3721: crom <= 108'o3722_3771_0006_4354_4007_0700_0000_0000_0000;
            12'o3722: crom <= 108'o3723_3333_0006_7174_4007_0700_0400_0000_0210;
            12'o3723: crom <= 108'o1060_3333_0004_7174_4007_0370_0400_0000_0212;
            12'o3724: crom <= 108'o3725_3333_0006_7174_4007_0700_0400_0000_0160;
            12'o3725: crom <= 108'o3726_3333_0006_7174_4007_0700_0400_0000_0161;
            12'o3726: crom <= 108'o1501_4571_1206_4374_4007_0700_0000_0036_0000;
            12'o3727: crom <= 108'o3730_4223_0000_4364_4277_0700_0200_0000_0010;
            12'o3730: crom <= 108'o3731_3551_1313_4374_0007_0700_0000_0002_4000;
            12'o3731: crom <= 108'o2532_4553_0600_4374_4007_0321_0000_0002_0000;
            12'o3732: crom <= 108'o3733_6551_0606_4374_0007_0700_0000_0000_1000;
            12'o3733: crom <= 108'o2534_3441_0605_4174_4007_0700_2000_0071_0007;
            12'o3734: crom <= 108'o2536_4553_1000_4374_4007_0321_0000_0000_0040;
            12'o3735: crom <= 108'o3736_3443_0300_4174_4007_0700_0200_0024_1016;
            12'o3736: crom <= 108'o1000_3771_0003_4365_5007_0700_0200_0000_0002;
            12'o3737: crom <= 108'o2572_4553_1300_4374_4007_0321_0000_0002_0000;
            12'o3740: crom <= 108'o2061_3771_0004_1276_6007_0701_0000_0000_1443;
            12'o3741: crom <= 108'o3456_0111_0703_4170_4007_0700_0210_0004_0012;
            12'o3742: crom <= 108'o3325_4571_1203_4374_4007_0700_0000_0077_7777;
            12'o3743: crom <= 108'o2156_3771_0006_1276_6007_0351_0000_0000_1443;
            12'o3744: crom <= 108'o3456_0111_0703_4174_4007_0700_0210_0004_0012;
            12'o3745: crom <= 108'o2576_4553_0600_4374_4007_0321_0000_0001_0000;
            12'o3746: crom <= 108'o3747_4221_0013_4170_4007_0700_0000_0000_0000;
            12'o3747: crom <= 108'o3750_3551_0606_4374_0007_0700_0000_0010_0000;
            12'o3750: crom <= 108'o2614_4553_1300_4374_4007_0321_0000_0000_4000;
            12'o3751: crom <= 108'o2111_3771_0006_0276_6007_0700_0000_0000_0000;
            12'o3752: crom <= 108'o1500_3111_0603_4174_4003_7700_0200_0003_0001;
            12'o3753: crom <= 108'o3755_3441_0305_4174_4007_0700_0000_0000_0000;
            12'o3754: crom <= 108'o2060_3771_0005_1276_6007_0701_0000_0000_1443;
            12'o3755: crom <= 108'o3756_5551_0305_4374_0007_0700_0000_0007_0000;
            12'o3756: crom <= 108'o3757_3443_0500_4174_4007_0701_0200_0000_0030;
            12'o3757: crom <= 108'o3760_4251_0404_4374_4007_0700_0000_0000_3777;
            12'o3760: crom <= 108'o3761_3551_0406_4374_4007_0700_0000_0040_0000;
            12'o3761: crom <= 108'o2616_4553_1300_4374_4007_0321_0000_0002_0000;
            12'o3762: crom <= 108'o3763_3771_0004_7274_4007_0701_0000_0000_0212;
            12'o3763: crom <= 108'o3764_3771_0005_7274_4007_0701_0000_0000_0213;
            12'o3764: crom <= 108'o3765_3771_0006_7274_4007_0701_0000_0000_0214;
            12'o3765: crom <= 108'o3766_3443_0300_4174_4007_0701_0200_0000_0032;
            12'o3766: crom <= 108'o0000_3771_0003_7274_4004_1701_0000_0000_0211;
            12'o3767: crom <= 108'o3770_3551_0304_4374_4007_0700_0000_0075_3777;
            12'o3770: crom <= 108'o3771_4111_0413_4174_0007_0700_0000_0000_0000;
            12'o3771: crom <= 108'o2630_3333_0003_4174_4007_0520_0000_0000_0000;
            12'o3772: crom <= 108'o2640_3443_0300_4174_4007_0370_0200_0024_1016;
            12'o3773: crom <= 108'o2644_4553_0300_4374_4007_0321_0000_0002_4000;
            12'o3774: crom <= 108'o2646_3333_0006_4174_4007_0520_0000_0000_0000;
            12'o3775: crom <= 108'o3776_3771_0004_4365_5007_0700_0200_0000_0002;
            12'o3776: crom <= 108'o2654_4553_0500_4374_4007_0331_0000_0000_0001;
            12'o3777: crom <= 108'o3720_3333_0003_7174_4007_0700_0400_0000_0211;
          endcase 
     end
endmodule
